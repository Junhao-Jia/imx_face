// Verilog netlist created by Tang Dynasty v6.0.135568
// Mon Jun  9 13:34:21 2025

`timescale 1ns / 1ps
module divider
  (
  clk,
  denominator,
  numerator,
  rst,
  start,
  done,
  quotient,
  remainder
  );

  input clk;
  input [31:0] denominator;
  input [47:0] numerator;
  input rst;
  input start;
  output done;
  output [47:0] quotient;
  output [31:0] remainder;

  parameter PIPLE = 50;
  parameter S_DEN = "UNSIGNED";
  parameter S_NUM = "UNSIGNED";
  parameter W_DEN = 32;
  parameter W_NUM = 48;
  parameter W_REM = 32;
  // localparam INPUT_PIPLINE = 1'b1;
  // localparam ITERA_PIPLINE = 48'b111111111111111111111111111111111111111111111111;
  // localparam OUTPUT_PIPLINE = 1'b1;
  // localparam SubSft[0].i = 0;
  // localparam SubSft[10].i = 10;
  // localparam SubSft[11].i = 11;
  // localparam SubSft[12].i = 12;
  // localparam SubSft[13].i = 13;
  // localparam SubSft[14].i = 14;
  // localparam SubSft[15].i = 15;
  // localparam SubSft[16].i = 16;
  // localparam SubSft[17].i = 17;
  // localparam SubSft[18].i = 18;
  // localparam SubSft[19].i = 19;
  // localparam SubSft[1].i = 1;
  // localparam SubSft[20].i = 20;
  // localparam SubSft[21].i = 21;
  // localparam SubSft[22].i = 22;
  // localparam SubSft[23].i = 23;
  // localparam SubSft[24].i = 24;
  // localparam SubSft[25].i = 25;
  // localparam SubSft[26].i = 26;
  // localparam SubSft[27].i = 27;
  // localparam SubSft[28].i = 28;
  // localparam SubSft[29].i = 29;
  // localparam SubSft[2].i = 2;
  // localparam SubSft[30].i = 30;
  // localparam SubSft[31].i = 31;
  // localparam SubSft[32].i = 32;
  // localparam SubSft[33].i = 33;
  // localparam SubSft[34].i = 34;
  // localparam SubSft[35].i = 35;
  // localparam SubSft[36].i = 36;
  // localparam SubSft[37].i = 37;
  // localparam SubSft[38].i = 38;
  // localparam SubSft[39].i = 39;
  // localparam SubSft[3].i = 3;
  // localparam SubSft[40].i = 40;
  // localparam SubSft[41].i = 41;
  // localparam SubSft[42].i = 42;
  // localparam SubSft[43].i = 43;
  // localparam SubSft[44].i = 44;
  // localparam SubSft[45].i = 45;
  // localparam SubSft[46].i = 46;
  // localparam SubSft[47].i = 47;
  // localparam SubSft[4].i = 4;
  // localparam SubSft[5].i = 5;
  // localparam SubSft[6].i = 6;
  // localparam SubSft[7].i = 7;
  // localparam SubSft[8].i = 8;
  // localparam SubSft[9].i = 9;
  wire [47:0] al_d3fd7d5a;
  wire [2:0] al_4b6a4daa;
  wire [68:0] al_6f9059d1;
  wire [47:0] al_f2b51288;
  wire [11:0] al_6a5d599;
  wire [47:0] al_5d497694;
  wire [10:0] al_fac191b8;
  wire [2:0] al_adb04807;
  wire [67:0] al_177a13cd;
  wire [47:0] al_6c6869d7;
  wire [12:0] al_2e720a5a;
  wire [47:0] al_c2901510;
  wire [11:0] al_c9ed4b28;
  wire [2:0] al_2e1bd9dc;
  wire [66:0] al_a6f4a789;
  wire [47:0] al_13d2e70f;
  wire [13:0] al_158480cc;
  wire [47:0] al_fb9cdc0e;
  wire [12:0] al_8fc8d46f;
  wire [2:0] al_c6d10c98;
  wire [65:0] al_515b933;
  wire [47:0] al_7cada4c1;
  wire [14:0] al_4f616992;
  wire [47:0] al_28d525d8;
  wire [13:0] al_a63aa325;
  wire [2:0] al_599810dd;
  wire [64:0] al_82ca84f8;
  wire [47:0] al_5fd65077;
  wire [15:0] al_e67d7d00;
  wire [47:0] al_8d341179;
  wire [14:0] al_1898703d;
  wire [2:0] al_903e8807;
  wire [63:0] al_297c219f;
  wire [47:0] al_174c5039;
  wire [16:0] al_e6544b06;
  wire [47:0] al_45052583;
  wire [15:0] al_ebfa785c;
  wire [2:0] al_5ed5f44b;
  wire [62:0] al_2e95330c;
  wire [47:0] al_1276f4f7;
  wire [17:0] al_eab6bdfe;
  wire [47:0] al_b5df9b8a;
  wire [16:0] al_b4daf6f3;
  wire [2:0] al_54284e1f;
  wire [61:0] al_b4e2b23b;
  wire [47:0] al_3692f86e;
  wire [18:0] al_7bf458d0;
  wire [47:0] al_28955387;
  wire [17:0] al_9c94ca47;
  wire [2:0] al_f83a6cd4;
  wire [60:0] al_e7d838f;
  wire [47:0] al_368cfa5b;
  wire [19:0] al_402e9e3e;
  wire [47:0] al_e55e130b;
  wire [18:0] al_def6d145;
  wire [2:0] al_b0a2efb7;
  wire [59:0] al_30e951fe;
  wire [47:0] al_e240f99f;
  wire [20:0] al_c49873a4;
  wire [47:0] al_abd7cd63;
  wire [19:0] al_bf1e6610;
  wire [2:0] al_3da4ff6f;
  wire [77:0] al_3bd314e4;
  wire [47:0] al_83a08f3f;
  wire [47:0] al_89f2771a;
  wire [1:0] al_33c3313d;
  wire [2:0] al_1c8da1e8;
  wire [58:0] al_e803eabe;
  wire [47:0] al_80a0f09e;
  wire [21:0] al_b2ee1d57;
  wire [47:0] al_cdad9264;
  wire [20:0] al_bd7f7f17;
  wire [2:0] al_acb3303d;
  wire [57:0] al_753f5f88;
  wire [47:0] al_98494645;
  wire [22:0] al_3e64f540;
  wire [47:0] al_f7ed724c;
  wire [21:0] al_be8c4478;
  wire [2:0] al_14a1a59a;
  wire [56:0] al_35594bd9;
  wire [47:0] al_bf34d64d;
  wire [23:0] al_365f90b4;
  wire [47:0] al_96533024;
  wire [22:0] al_f1d740ba;
  wire [2:0] al_21143207;
  wire [55:0] al_f2bb4ec4;
  wire [47:0] al_f0f43754;
  wire [24:0] al_21ee8bc;
  wire [47:0] al_e60d8647;
  wire [23:0] al_d3734717;
  wire [2:0] al_e0dc7e9e;
  wire [54:0] al_3029c49a;
  wire [47:0] al_86280a69;
  wire [25:0] al_511419f7;
  wire [47:0] al_f78b30ce;
  wire [24:0] al_4a4fb8f1;
  wire [2:0] al_bade9fae;
  wire [53:0] al_5181785e;
  wire [47:0] al_9e3033a4;
  wire [26:0] al_693e712c;
  wire [47:0] al_63579c4c;
  wire [25:0] al_28f9bf01;
  wire [2:0] al_8f9ab06;
  wire [52:0] al_6a56028d;
  wire [47:0] al_7397600a;
  wire [27:0] al_cabe3087;
  wire [47:0] al_2c297489;
  wire [26:0] al_c0ef3ebf;
  wire [2:0] al_fee4bd37;
  wire [51:0] al_b6768e55;
  wire [47:0] al_e4be4089;
  wire [28:0] al_c307e46;
  wire [47:0] al_9857f6b5;
  wire [27:0] al_d71a2aba;
  wire [2:0] al_e0e2aae4;
  wire [50:0] al_222a5f4d;
  wire [47:0] al_4a463b38;
  wire [29:0] al_794ac8f;
  wire [47:0] al_e343d659;
  wire [28:0] al_c7a3cd65;
  wire [2:0] al_5db428bb;
  wire [49:0] al_d1a07609;
  wire [47:0] al_32ba5b24;
  wire [30:0] al_af127331;
  wire [47:0] al_14165a56;
  wire [29:0] al_bad3f013;
  wire [2:0] al_67f5b0b3;
  wire [76:0] al_6a637a32;
  wire [47:0] al_3d0cfeb4;
  wire [47:0] al_a9b28455;
  wire [2:0] al_b54c1014;
  wire [2:0] al_8d805738;
  wire [48:0] al_627988c3;
  wire [47:0] al_690b21a4;
  wire [31:0] al_2c47200f;
  wire [47:0] al_3ccb3a4f;
  wire [30:0] al_9d67405f;
  wire [2:0] al_74993dd2;
  wire [47:0] al_a5e9c08d;
  wire [47:0] al_57dc9b0c;
  wire [32:0] al_d8106c92;
  wire [47:0] al_eb7d14b9;
  wire [31:0] al_b40233aa;
  wire [2:0] al_2e2a074f;
  wire [46:0] al_930eb7ed;
  wire [47:0] al_e7fdd367;
  wire [33:0] al_ede1be73;
  wire [47:0] al_f100da9b;
  wire [32:0] al_586198c7;
  wire [2:0] al_ad601da1;
  wire [45:0] al_400c3c08;
  wire [46:0] al_5675a322;
  wire [33:0] al_2232b9e8;
  wire [46:0] al_dacf1710;
  wire [33:0] al_3a0a3044;
  wire [2:0] al_ff0af5c2;
  wire [44:0] al_304b2866;
  wire [45:0] al_c7be2582;
  wire [33:0] al_fab6b65e;
  wire [45:0] al_be68a6d4;
  wire [34:0] al_64e3fb17;
  wire [2:0] al_65c09044;
  wire [43:0] al_bac230e2;
  wire [44:0] al_d99b0302;
  wire [33:0] al_cc14d64d;
  wire [44:0] al_b75cf8f9;
  wire [35:0] al_8642d51e;
  wire [2:0] al_4c0a9e6a;
  wire [42:0] al_ccda870f;
  wire [43:0] al_cb972596;
  wire [33:0] al_35eab049;
  wire [43:0] al_dd187023;
  wire [36:0] al_29052500;
  wire [2:0] al_88b72b17;
  wire [41:0] al_8c4c0e00;
  wire [42:0] al_7848278f;
  wire [33:0] al_c73a14b6;
  wire [42:0] al_b8e7a164;
  wire [37:0] al_6cd22c9c;
  wire [2:0] al_d72cf58c;
  wire [40:0] al_a32146c7;
  wire [41:0] al_ab78d0a0;
  wire [33:0] al_d4021fa0;
  wire [41:0] al_1dac5d46;
  wire [38:0] al_5dd36af2;
  wire [2:0] al_90e1f6ef;
  wire [39:0] al_2ecc3265;
  wire [40:0] al_7af0d249;
  wire [33:0] al_1d982a67;
  wire [40:0] al_d9c08430;
  wire [39:0] al_b6775e93;
  wire [2:0] al_44882eca;
  wire [75:0] al_b052c226;
  wire [47:0] al_592f1b09;
  wire [47:0] al_8c015879;
  wire [3:0] al_b18b7cbb;
  wire [2:0] al_5bcbf559;
  wire [38:0] al_615b2119;
  wire [39:0] al_ce3b275;
  wire [33:0] al_79977513;
  wire [39:0] al_92415709;
  wire [40:0] al_56efbba9;
  wire [2:0] al_16eefd24;
  wire [37:0] al_aa3e519e;
  wire [38:0] al_f8daefdd;
  wire [33:0] al_a972f2b7;
  wire [38:0] al_c5d46f6b;
  wire [41:0] al_3357c8f6;
  wire [2:0] al_993138f9;
  wire [36:0] al_5e4a13f0;
  wire [37:0] al_32798732;
  wire [33:0] al_a7bae927;
  wire [37:0] al_93803eaa;
  wire [42:0] al_7d914746;
  wire [2:0] al_d5d72c9e;
  wire [35:0] al_22838ccb;
  wire [36:0] al_2f60c4e5;
  wire [33:0] al_6c10dd8f;
  wire [36:0] al_1a0e1c89;
  wire [43:0] al_97fb94a7;
  wire [2:0] al_2be1e26f;
  wire [34:0] al_44122f34;
  wire [35:0] al_167f3ebe;
  wire [33:0] al_a352434c;
  wire [35:0] al_7452903f;
  wire [44:0] al_c2cdf2f1;
  wire [2:0] al_5d2b923b;
  wire [33:0] al_7e0865ed;
  wire [34:0] al_cafe0ad;
  wire [33:0] al_fc56973;
  wire [34:0] al_ce2f96cc;
  wire [45:0] al_2c312a8;
  wire [2:0] al_1fd6d456;
  wire [32:0] al_8ee40da8;
  wire [33:0] al_13d036ce;
  wire [33:0] al_65caf2b5;
  wire [33:0] al_b328a515;
  wire [46:0] al_f3197cbe;
  wire [2:0] al_7a934789;
  wire [31:0] al_ac1cba4d;
  wire [32:0] al_8f041238;
  wire [32:0] al_4101ed12;
  wire [33:0] al_42247ac7;
  wire [47:0] al_59124752;
  wire [2:0] al_f336c405;
  wire [74:0] al_28202fa7;
  wire [47:0] al_1d4399b1;
  wire [47:0] al_7a8c14f1;
  wire [4:0] al_917df14b;
  wire [2:0] al_f23786d8;
  wire [73:0] al_68bb3ebd;
  wire [47:0] al_1b3e91c5;
  wire [6:0] al_504aeee4;
  wire [47:0] al_7d7cdb8e;
  wire [5:0] al_4682e2e2;
  wire [2:0] al_6e4d5f5f;
  wire [72:0] al_f2a9de02;
  wire [47:0] al_15503509;
  wire [7:0] al_b9ac5fd4;
  wire [47:0] al_78306f09;
  wire [6:0] al_22a22ff3;
  wire [2:0] al_d255f877;
  wire [71:0] al_5206392b;
  wire [47:0] al_59bef53b;
  wire [8:0] al_f87eab88;
  wire [47:0] al_601b9c02;
  wire [7:0] al_9c3e2402;
  wire [2:0] al_30922aac;
  wire [70:0] al_d6cb04b6;
  wire [47:0] al_f7a9a92b;
  wire [9:0] al_5b8748c3;
  wire [47:0] al_3b7f0416;
  wire [8:0] al_4dd3fb65;
  wire [2:0] al_36d845bb;
  wire [69:0] al_c1960abd;
  wire [47:0] al_5283b07c;
  wire [10:0] al_93772c3;
  wire [47:0] al_bcaebe78;
  wire [9:0] al_3cd0a9ea;
  wire [2:0] al_dc871c53;
  wire [78:0] al_9d1d5c0;
  wire [47:0] al_a5806bc7;
  wire [47:0] al_bfaf4e7;
  wire [47:0] al_3b63a678;
  wire al_51794c84;
  wire al_147773d6;
  wire al_56e18a80;
  wire al_1435a49e;
  wire al_e0cc30a4;
  wire al_1e3141cc;
  wire al_4a4b505;
  wire al_e8aefc81;
  wire al_689ce8c2;
  wire al_b32218f4;
  wire al_aa787729;
  wire al_c9b85978;
  wire al_1472bf2f;
  wire al_787b0a64;
  wire al_c3020830;
  wire al_fa8bcfd;
  wire al_258d6ce0;
  wire al_dc10836c;
  wire al_4de5b5ba;
  wire al_1a08a0b7;
  wire al_fe80d5e5;
  wire al_56ca40b1;
  wire al_2f2f061f;
  wire al_75e67c73;
  wire al_93654000;
  wire al_95c9121c;
  wire al_6a7cf4f6;
  wire al_7d43f9f9;
  wire al_c2244c00;
  wire al_3690d0d4;
  wire al_5b92a62d;
  wire al_59478e92;
  wire al_9ea91fcd;
  wire al_3d9987d2;
  wire al_c5d02c43;
  wire al_8889fefd;
  wire al_28b0e45b;
  wire al_1e2e550f;
  wire al_3afa0b96;
  wire al_c029c247;
  wire al_62aba81a;
  wire al_e889058f;
  wire al_82230b41;
  wire al_88df3967;
  wire al_2824b693;
  wire al_6d794600;
  wire al_6e4bbf49;
  wire al_2ef9708;
  wire al_f452a7c;
  wire al_32e1725d;
  wire al_a83c9088;
  wire al_f9a74458;
  wire al_54803b10;
  wire al_7ba0f244;
  wire al_4e9b63c9;
  wire al_dcea9b4;
  wire al_afad458d;
  wire al_90e336e1;
  wire al_d41ac52e;
  wire al_2bfcf033;
  wire al_bf8f4b75;
  wire al_98398e18;
  wire al_463946df;
  wire al_967a5f00;
  wire al_110841cf;
  wire al_9bebb94b;
  wire al_e2402cc4;
  wire al_49617358;
  wire al_f9d08351;
  wire al_57db75f0;
  wire al_b261805d;
  wire al_d2377beb;
  wire al_f58e7482;
  wire al_2576177;
  wire al_64c2879;
  wire al_6b5869dc;
  wire al_f6f2dce7;
  wire al_9cb945d3;
  wire al_c0342edb;
  wire al_abf1ad7c;
  wire al_3971206e;
  wire al_36535fd3;
  wire al_430e5cec;
  wire al_35bf8c77;
  wire al_6a165344;
  wire al_edeaa856;
  wire al_f3dfd21a;
  wire al_b398ed4f;
  wire al_5c1aec80;
  wire al_1c3eecd0;
  wire al_62e1f39;
  wire al_ee6cfa1b;
  wire al_7e84b0e7;
  wire al_36b609cf;
  wire al_e216e162;
  wire al_436534ab;
  wire al_1a52e2b9;
  wire al_1686893d;
  wire al_8c362b8c;
  wire al_ca0bc000;
  wire al_631fb54;
  wire al_6a2b173c;
  wire al_c111311e;
  wire al_a67d66f1;
  wire al_5cbcdb58;
  wire al_bb2c445c;
  wire al_a217d3f1;
  wire al_5cde9409;
  wire al_7b31c923;
  wire al_855bfb89;
  wire al_c41c8842;
  wire al_29e9ad49;
  wire al_786a64be;
  wire al_9b1b3762;
  wire al_371bfa10;
  wire al_eea0690a;
  wire al_670e1d07;
  wire al_ee69ef7a;
  wire al_11e5467d;
  wire al_3910e4e4;
  wire al_35b24b05;
  wire al_61d00fc7;
  wire al_550f60c3;
  wire al_5f55c3b4;
  wire al_dc7a89a9;
  wire al_5aec0d3d;
  wire al_146c9954;
  wire al_95294fb6;
  wire al_2b309dfb;
  wire al_af8062a0;
  wire al_3c2e3c3a;
  wire al_b4c76c23;
  wire al_bcaace37;
  wire al_6dbf3665;
  wire al_8a54e775;
  wire al_8f1f7251;
  wire al_eb782a2a;
  wire al_d3a3aa84;
  wire al_43acb4d3;
  wire al_2a00900c;
  wire al_66810f7a;
  wire al_dbcf415b;
  wire al_e40ec610;
  wire al_3ca88873;
  wire al_4ff8e4;
  wire al_cd79137f;
  wire al_dbca7fa0;
  wire al_547f2817;
  wire al_85dc8a57;
  wire al_2ed9b6e7;
  wire al_283f9817;
  wire al_1967a37e;
  wire al_32707238;
  wire al_2c79b8f0;
  wire al_6fa79631;
  wire al_683a8463;
  wire al_c6efb15f;
  wire al_16cee9f7;
  wire al_33147ecd;
  wire al_7644ebe6;
  wire al_a21a5b9f;
  wire al_84143d7e;
  wire al_2e9e4aac;
  wire al_a7eb7389;
  wire al_122ce731;
  wire al_93a235f1;
  wire al_bfc9143c;
  wire al_8e30be98;
  wire al_2ee33b11;
  wire al_cc4f6241;
  wire al_27369a88;
  wire al_790961ba;
  wire al_ed8719fc;
  wire al_21a14027;
  wire al_f719f95a;
  wire al_eb9006e0;
  wire al_6680c576;
  wire al_7820cd3f;
  wire al_91e67405;
  wire al_1f539415;
  wire al_fdf27789;
  wire al_cd1eb597;
  wire al_95c541ba;
  wire al_c62ed6f3;
  wire al_2e458e8c;
  wire al_314816f3;
  wire al_3db819db;
  wire al_4cb58e58;
  wire al_61f7300c;
  wire al_51cbf969;
  wire al_31d377e1;
  wire al_5e3c7f1a;
  wire al_67c30993;
  wire al_1c99d5f6;
  wire al_66df73c7;
  wire al_a3e63ee7;
  wire al_63d267c1;
  wire al_8aa456b9;
  wire al_7fa59108;
  wire al_54c1a264;
  wire al_1937c3b1;
  wire al_8d689511;
  wire al_24deb4a;
  wire al_38e8d651;
  wire al_456aad79;
  wire al_26b2c4d9;
  wire al_9780212c;
  wire al_93d510f7;
  wire al_7cbeb255;
  wire al_5303c8c4;
  wire al_e8916352;
  wire al_1634b160;
  wire al_2d07102b;
  wire al_3b0f07fc;
  wire al_45fda30c;
  wire al_ca8a5a31;
  wire al_fd5ea84d;
  wire al_ff28a985;
  wire al_b8462556;
  wire al_54775a2b;
  wire al_39d57d97;
  wire al_e98f3c34;
  wire al_5761f230;
  wire al_2283cfcc;
  wire al_5d7328e8;
  wire al_93496304;
  wire al_abc34969;
  wire al_90929116;
  wire al_2da51efc;
  wire al_c89089ad;
  wire al_e37f1d18;
  wire al_77a0ba2a;
  wire al_c1b434db;
  wire al_5622df9b;
  wire al_e3ce0c99;
  wire al_7a39fd90;
  wire al_290a897c;
  wire al_39495ba2;
  wire al_ff8767e1;
  wire al_edbcd561;
  wire al_b68658c6;
  wire al_7bc5cf46;
  wire al_c9c0b8e5;
  wire al_ddf57730;
  wire al_bcf04c60;
  wire al_76e6b917;
  wire al_f66e0990;
  wire al_c0b6cd6e;
  wire al_5507d757;
  wire al_216ce40;
  wire al_66aff298;
  wire al_cdeed011;
  wire al_d2fa64e6;
  wire al_e0707d5b;
  wire al_b9091bb4;
  wire al_cafa3568;
  wire al_177f9d69;
  wire al_8d529875;
  wire al_663d37b6;
  wire al_bd5caa9f;
  wire al_95b12900;
  wire al_a9d8f8;
  wire al_3459937f;
  wire al_b062dbda;
  wire al_ab1c35b3;
  wire al_41371141;
  wire al_a7492340;
  wire al_8f25dca0;
  wire al_b27b3769;
  wire al_a8fb6998;
  wire al_18a0a383;
  wire al_2f3a1692;
  wire al_d4bc7f3e;
  wire al_72d62b1c;
  wire al_4e56a0da;
  wire al_1240f9a6;
  wire al_2ec3de14;
  wire al_b48c402a;
  wire al_63f814e;
  wire al_3c4a2199;
  wire al_f832136c;
  wire al_934e501;
  wire al_d460c819;
  wire al_88e1bda3;
  wire al_1821d93d;
  wire al_b4ee9e86;
  wire al_9828f0b3;
  wire al_3f6c8445;
  wire al_28e359b1;
  wire al_4b337999;
  wire al_92297df8;
  wire al_7dcd3618;
  wire al_68deb8d6;
  wire al_274f6baa;
  wire al_86dc2d65;
  wire al_f4230bb8;
  wire al_ada1b083;
  wire al_5051b702;
  wire al_fd100c07;
  wire al_f492d664;
  wire al_6d3aa56f;
  wire al_534497b1;
  wire al_cb73325b;
  wire al_b65c9b4;
  wire al_178c71f6;
  wire al_cbbef4f;
  wire al_9e9b738f;
  wire al_a076256b;
  wire al_7930e629;
  wire al_a521f9f;
  wire al_5f29b438;
  wire al_3ce4b2fd;
  wire al_86766b99;
  wire al_b17e5f2d;
  wire al_a2b56c4c;
  wire al_998abf81;
  wire al_ce61dd12;
  wire al_1ae1e567;
  wire al_eea1c0b5;
  wire al_8d1ae89a;
  wire al_92faecea;
  wire al_ddf49d7d;
  wire al_5613036;
  wire al_c86a97ab;
  wire al_ac57c034;
  wire al_920c4e9a;
  wire al_1283ff0b;
  wire al_44359cb4;
  wire al_1fc8de48;
  wire al_9b620d8d;
  wire al_c5542b59;
  wire al_fef84737;
  wire al_d8cfcc23;
  wire al_96385301;
  wire al_2021f859;
  wire al_86a4ed5a;
  wire al_52f700f5;
  wire al_1024eced;
  wire al_55cc2fd4;
  wire al_58146106;
  wire al_b0f0b903;
  wire al_f01ea45c;
  wire al_2b0b3830;
  wire al_cc9bf94;
  wire al_4a3ef4b7;
  wire al_168ee139;
  wire al_c52a2c84;
  wire al_3a745b61;
  wire al_328e2c2d;
  wire al_86e77cd0;
  wire al_8b31527f;
  wire al_1119be30;
  wire al_71939d74;
  wire al_d3344326;
  wire al_e466bfff;
  wire al_fe06d9ee;
  wire al_79cadb17;
  wire al_e2799097;
  wire al_12391d73;
  wire al_e4135f97;
  wire al_7c91f33c;
  wire al_5576ac23;
  wire al_3f791172;
  wire al_1c1093cd;
  wire al_61436e1a;
  wire al_bedba12b;
  wire al_c3463f35;
  wire al_fa3d49c2;
  wire al_caf86cb;
  wire al_603373a4;
  wire al_236d63a;
  wire al_1e576ba8;
  wire al_79f81494;
  wire al_921bd39c;
  wire al_38de2714;
  wire al_b7b5bdbe;
  wire al_d7aedbc5;
  wire al_43e60c58;
  wire al_f67fc030;
  wire al_e1b1f9c7;
  wire al_d27a6f7e;
  wire al_7932b374;
  wire al_93343d44;
  wire al_563f66f8;
  wire al_eb1ae9e7;
  wire al_e483a091;
  wire al_c3dfa0bb;
  wire al_f67f9b7;
  wire al_a6e65c64;
  wire al_a7b28424;
  wire al_17c9f81e;
  wire al_ff089b0;
  wire al_7f19c0cd;
  wire al_aadee294;
  wire al_1f32676d;
  wire al_e995362;
  wire al_28383266;
  wire al_d33bf669;
  wire al_c70e8ffd;
  wire al_f531391e;
  wire al_c1cd2e91;
  wire al_5361b136;
  wire al_1f83c861;
  wire al_1fd9ea3c;
  wire al_e10dc145;
  wire al_dec1a002;
  wire al_9e36993d;
  wire al_8302a2a2;
  wire al_78579729;
  wire al_cce3e61c;
  wire al_edfe5545;
  wire al_8afadf84;
  wire al_91c4f866;
  wire al_dfb38e7;
  wire al_ea5a8045;
  wire al_5594316d;
  wire al_802edd1b;
  wire al_4ed141e3;
  wire al_a9bde1cf;
  wire al_b879dc6c;
  wire al_8f601d11;
  wire al_1861ccb9;
  wire al_417b1b7f;
  wire al_a4400d46;
  wire al_59eab12e;
  wire al_1af64e4d;
  wire al_ecd39a7;
  wire al_a7d6fdcd;
  wire al_7de07321;
  wire al_df148873;
  wire al_1f49b9e4;
  wire al_832fb3e;
  wire al_2d137dff;
  wire al_fd484a6d;
  wire al_1d7722f2;
  wire al_83dc3e4f;
  wire al_e7c4a377;
  wire al_153001b0;
  wire al_90b73cc5;
  wire al_6cc49207;
  wire al_88ebd806;
  wire al_9ba3e8a0;
  wire al_c1436409;
  wire al_a907358b;
  wire al_7c92a6e7;
  wire al_2848275b;
  wire al_1cb31d61;
  wire al_ddf9bf5e;
  wire al_4cef4276;
  wire al_6cf3b362;
  wire al_e0b0ba1d;
  wire al_5c52a055;
  wire al_90d0cde9;
  wire al_b506c4;
  wire al_63ccb9ff;
  wire al_72ec7913;
  wire al_a727e78e;
  wire al_61742d3d;
  wire al_da23077d;
  wire al_d907d72;
  wire al_941ec574;
  wire al_e915b010;
  wire al_4f44504e;
  wire al_30d605ba;
  wire al_8c151872;
  wire al_e2a656fd;
  wire al_55ab11c1;
  wire al_281a7b5c;
  wire al_17661190;
  wire al_ba73d945;
  wire al_7e55c045;
  wire al_efd0595d;
  wire al_83ddd85b;
  wire al_4697075e;
  wire al_5ad7048f;
  wire al_9071f0e5;
  wire al_e5398263;
  wire al_b191d1e0;
  wire al_49a0e61d;
  wire al_86984010;
  wire al_862cc7f8;
  wire al_b980f13c;
  wire al_db4a0b3b;
  wire al_b7c44457;
  wire al_c68c13d2;
  wire al_f144ba04;
  wire al_2e50ac1e;
  wire al_e418756e;
  wire al_8653cc11;
  wire al_fa5db848;
  wire al_39ade860;
  wire al_7183147;
  wire al_616fbe10;
  wire al_47d76c66;
  wire al_ebfbc5f1;
  wire al_3f596b4e;
  wire al_4b8b49e0;
  wire al_608458c0;
  wire al_14b22db9;
  wire al_f04c5c1a;
  wire al_6b3dc9d;
  wire al_b33cc591;
  wire al_b34ec3bf;
  wire al_eb58c5cb;
  wire al_95542881;
  wire al_8b31dee3;
  wire al_1c1f1cb1;
  wire al_55f734a7;
  wire al_51e8603;
  wire al_ffbd9e7e;
  wire al_2aef1337;
  wire al_a3fc3ebc;
  wire al_5cdd85d5;
  wire al_1add508;
  wire al_5a84d22c;
  wire al_cf720ce3;
  wire al_656d5c84;
  wire al_de32c090;
  wire al_f42fa6ce;
  wire al_b6af5571;
  wire al_c2ee5e5b;
  wire al_43f00cc1;
  wire al_a541ec8a;
  wire al_74501eb3;
  wire al_ffc5f376;
  wire al_d3b64099;
  wire al_9abafd70;
  wire al_8225507c;
  wire al_ff92482;
  wire al_2e13f976;
  wire al_bd65eabf;
  wire al_ede5673b;
  wire al_70a9c221;
  wire al_532cc9a8;
  wire al_ea82bb3a;
  wire al_d637b77b;
  wire al_2e7f5ba5;
  wire al_93b7a367;
  wire al_3d8d5fa3;
  wire al_294cc864;
  wire al_3220468;
  wire al_b1e53313;
  wire al_e4e8fccd;
  wire al_d45bda05;
  wire al_50a889e9;
  wire al_45125ed0;
  wire al_256e1d30;
  wire al_6b8e1d26;
  wire al_b57afe80;
  wire al_34a605a;
  wire al_56bd060e;
  wire al_c328a853;
  wire al_4ffec454;
  wire al_d37de394;
  wire al_1b2a14dc;
  wire al_31a7b4b6;
  wire al_d2a76de7;
  wire al_53f78588;
  wire al_89b70b3b;
  wire al_15cd8a93;
  wire al_eb481677;
  wire al_1b3445fd;
  wire al_1ab93794;
  wire al_c1f5ea1e;
  wire al_57899523;
  wire al_94297415;
  wire al_1f080dc4;
  wire al_de10dc85;
  wire al_b42d0d53;
  wire al_fd6c2091;
  wire al_c10da5dd;
  wire al_dd5f2a54;
  wire al_11eefeb5;
  wire al_64eb948d;
  wire al_6ed7702d;
  wire al_f68e810e;
  wire al_430afd8b;
  wire al_f0ecaeb6;
  wire al_1376bcb0;
  wire al_4a06e815;
  wire al_58a18b68;
  wire al_4085a271;
  wire al_858f1c0c;
  wire al_364abc0a;
  wire al_9909f3ca;
  wire al_bacdad1b;
  wire al_9bec1f33;
  wire al_83f595b;
  wire al_91824dca;
  wire al_9ba07719;
  wire al_fc839793;
  wire al_739af9ca;
  wire al_de14f218;
  wire al_112db54d;
  wire al_f31a4cd8;
  wire al_a77da9ed;
  wire al_9d63b53d;
  wire al_b187ff7c;
  wire al_a416feb9;
  wire al_3a2fee85;
  wire al_af90c070;
  wire al_a9f17098;
  wire al_7b8d96e2;
  wire al_a5b3371d;
  wire al_aa3a575d;
  wire al_354eea5a;
  wire al_94b0c7d1;
  wire al_cbca04a4;
  wire al_9767aad8;
  wire al_1fe3c2d1;
  wire al_b233479;
  wire al_71be4cd6;
  wire al_54a79559;
  wire al_c4782520;
  wire al_b1f716e3;
  wire al_a59de26c;
  wire al_561ce4c4;
  wire al_2451e527;
  wire al_2bed1d6f;
  wire al_a9898f67;
  wire al_7999a920;
  wire al_dcd3196f;
  wire al_9d1db55;
  wire al_9240c8a4;
  wire al_f5953bb1;
  wire al_ff96e0f;
  wire al_fdc157ff;
  wire al_fa3f4f58;
  wire al_f0643c82;
  wire al_1106f695;
  wire al_474d64a7;
  wire al_d079fcc4;
  wire al_8af08334;
  wire al_d3786c88;
  wire al_1c2d1a70;
  wire al_47dadb08;
  wire al_4145de8a;
  wire al_1dddd2e5;
  wire al_90ad6b5d;
  wire al_f4e9ff5b;
  wire al_615d34bc;
  wire al_7b56c629;
  wire al_90865e32;
  wire al_5bc29d76;
  wire al_b89115b;
  wire al_1bed3aa5;
  wire al_ee91a42b;
  wire al_d9039a1f;
  wire al_5dced79d;
  wire al_c2c29ff3;
  wire al_bb679170;
  wire al_e9214bad;
  wire al_a13e1232;
  wire al_e9639971;
  wire al_15e685d4;
  wire al_d09dedfa;
  wire al_d38c342e;
  wire al_718df034;
  wire al_97f6d29;
  wire al_d87faa07;
  wire al_f45a16f4;
  wire al_23c32ed1;
  wire al_5c729632;
  wire al_117d184b;
  wire al_cd65094;
  wire al_cdc4fc2e;
  wire al_88c69413;
  wire al_624a5f2d;
  wire al_d71b24d6;
  wire al_a1d5dec3;
  wire al_12dadb42;
  wire al_bc1185ef;
  wire al_d5531fd2;
  wire al_b07fbb26;
  wire al_8a3c5223;
  wire al_4dd1780b;
  wire al_a06e1c18;
  wire al_50022df0;
  wire al_58ce9b0f;
  wire al_542e503f;
  wire al_55bbc798;
  wire al_aa5ae88a;
  wire al_5b4dd00b;
  wire al_584eea74;
  wire al_c6e57848;
  wire al_efc6812a;
  wire al_10825af9;
  wire al_bbfa0f21;
  wire al_bf9072a4;
  wire al_18cc4352;
  wire al_cd59a509;
  wire al_a9bd067e;
  wire al_8ff81b47;
  wire al_91d9bc15;
  wire al_da758300;
  wire al_44b995d2;
  wire al_f3c33aa1;
  wire al_1b86bf86;
  wire al_d1142aec;
  wire al_6600d0f4;
  wire al_e73d5abc;
  wire al_a2618249;
  wire al_e181fe09;
  wire al_c77349a0;
  wire al_f63d2d13;
  wire al_46537d2e;
  wire al_a889f4bf;
  wire al_accde4d;
  wire al_508bf5eb;
  wire al_e82cb205;
  wire al_4f99c2a2;
  wire al_46d116b1;
  wire al_7a5c8d6e;
  wire al_86d44bba;
  wire al_53b3d48f;
  wire al_7ed64a67;
  wire al_779d4335;
  wire al_e0b2aa1b;
  wire al_38a13889;
  wire al_8419f2ed;
  wire al_f54b9335;
  wire al_8ed6d91d;
  wire al_3a63fdce;
  wire al_7d6eed39;
  wire al_ebfc32c7;
  wire al_34381ac;
  wire al_49175cff;
  wire al_63ff6480;
  wire al_27dd2411;
  wire al_a911db93;
  wire al_405a9f2c;
  wire al_e8221400;
  wire al_a28a7cde;
  wire al_61046848;
  wire al_51208526;
  wire al_93c8ec69;
  wire al_52ebcad4;
  wire al_ed6494a;
  wire al_7d39bb7d;
  wire al_22aeb069;
  wire al_5d314c19;
  wire al_53a672a;
  wire al_39309161;
  wire al_9a288672;
  wire al_d2d28755;
  wire al_baeae313;
  wire al_63993f05;
  wire al_b24d98eb;
  wire al_89a36400;
  wire al_1a8ff40a;
  wire al_585d083c;
  wire al_bada19ee;
  wire al_3184f1ad;
  wire al_2bfc7bfc;
  wire al_e59a7f64;
  wire al_5a56dd8c;
  wire al_c8cc3a74;
  wire al_2a0ec313;
  wire al_e6e3c466;
  wire al_d781087a;
  wire al_8cba2b5a;
  wire al_cb8ad3a1;
  wire al_3c5da63;
  wire al_731d9b96;
  wire al_bf6ae1e2;
  wire al_714663e5;
  wire al_4cf28725;
  wire al_639c27a1;
  wire al_c465640a;
  wire al_d013c2db;
  wire al_86c1a1f7;
  wire al_e412eb65;
  wire al_f01a65dd;
  wire al_e6ba2112;
  wire al_3fdd05cb;
  wire al_43bdc053;
  wire al_be037ee1;
  wire al_e6e34f55;
  wire al_a638954c;
  wire al_9eeedd82;
  wire al_58c037cd;
  wire al_f841ecaa;
  wire al_e7643d65;
  wire al_d681bdcc;
  wire al_537d0180;
  wire al_c18839e1;
  wire al_a12bfe23;
  wire al_23bcebc4;
  wire al_94fa0ad9;
  wire al_3773fc04;
  wire al_8eedc273;
  wire al_bd0a1f9d;
  wire al_48931d43;
  wire al_bc9b0eaa;
  wire al_35d02980;
  wire al_fee10e00;
  wire al_56671d76;
  wire al_912d325d;
  wire al_9f5bba13;
  wire al_93b8640e;
  wire al_e3447775;
  wire al_ba94a953;
  wire al_75a96ab5;
  wire al_3c16a30a;
  wire al_fdf3ddc7;
  wire al_2c40a92e;
  wire al_d57289de;
  wire al_c0464485;
  wire al_6cd1bb56;
  wire al_805eafcd;
  wire al_afc2f09b;
  wire al_b626be09;
  wire al_47857556;
  wire al_cdf5386d;
  wire al_44a63fb7;
  wire al_d8fe84e6;
  wire al_6d9bce46;
  wire al_46c8a269;
  wire al_ba4595c0;
  wire al_5bf37252;
  wire al_8cb44011;
  wire al_b5df3e43;
  wire al_2392f558;
  wire al_7581bd0d;
  wire al_f01e9810;
  wire al_4b0822cb;
  wire al_46ca2999;
  wire al_f327e49f;
  wire al_6af99fb0;
  wire al_f9708799;
  wire al_ce755696;
  wire al_8ceeb1d6;
  wire al_56f936a;
  wire al_c17b3665;
  wire al_4942e686;
  wire al_fa0cd080;
  wire al_b938610a;
  wire al_76221ee1;
  wire al_73d542b1;
  wire al_a0e7f496;
  wire al_5516d10;
  wire al_cade3756;
  wire al_dc3daad0;
  wire al_cf98adbf;
  wire al_b30ebdf6;
  wire al_2258030e;
  wire al_8bfba661;
  wire al_9e4c11b8;
  wire al_7116cd2;
  wire al_7c2f83cb;
  wire al_689a4219;
  wire al_6d6bb647;
  wire al_d9a99e6d;
  wire al_d98a025f;
  wire al_6272599f;
  wire al_c512c49;
  wire al_40c30b4d;
  wire al_de3e7627;
  wire al_92ccaa05;
  wire al_40670ee4;
  wire al_12b84efd;
  wire al_7d13d94f;
  wire al_b458e911;
  wire al_f5397afe;
  wire al_626a930b;
  wire al_3bcfaff1;
  wire al_4059e403;
  wire al_ab96385b;
  wire al_b2787015;
  wire al_e23a271f;
  wire al_eed33fc3;
  wire al_7e086938;
  wire al_4ebf21a;
  wire al_f74ec05f;
  wire al_b1a4aa4;
  wire al_98dec4e;
  wire al_2825c36a;
  wire al_ca256ef5;
  wire al_cac22815;
  wire al_7b366c25;
  wire al_306af3cf;
  wire al_4957c6a5;
  wire al_8a47c612;
  wire al_f65c10;
  wire al_6a66d91e;
  wire al_bcbd4e1b;
  wire al_792f9fb1;
  wire al_1f9c650e;
  wire al_e88204f;
  wire al_c435b5e6;
  wire al_13c84cc8;
  wire al_21c2c54f;
  wire al_fe48089b;
  wire al_fe0b2c2e;
  wire al_8b619c3b;
  wire al_a522c3d4;
  wire al_e347376a;
  wire al_28f6cbc1;
  wire al_17617f0f;
  wire al_510c2901;
  wire al_8aca8bdd;
  wire al_94c5d51b;
  wire al_ec8c91da;
  wire al_a1bb6a32;
  wire al_ac09860;
  wire al_8818311f;
  wire al_189a7687;
  wire al_b94ff95a;
  wire al_1a56b969;
  wire al_5971bdb0;
  wire al_a1353883;
  wire al_a8675d43;
  wire al_2dcd8322;
  wire al_1e9d53ff;
  wire al_a3e2ac47;
  wire al_da3e5716;
  wire al_6b874685;
  wire al_ab74a1e3;
  wire al_6c10ec91;
  wire al_c829298;
  wire al_88013228;
  wire al_ebe24e3d;
  wire al_c22e023d;
  wire al_7aed21eb;
  wire al_de434a70;
  wire al_4026dc20;
  wire al_7c090755;
  wire al_ae7b2873;
  wire al_e8aded2c;
  wire al_d89660dd;
  wire al_a0eacc1c;
  wire al_371958b8;
  wire al_69ee2d7e;
  wire al_a313220b;
  wire al_cde03fa5;
  wire al_47e767;
  wire al_160b1ef;
  wire al_8178bce7;
  wire al_ebc6f995;
  wire al_bc6f54a9;
  wire al_1a110913;
  wire al_b4aada3d;
  wire al_5f7332b4;
  wire al_64d12b15;
  wire al_13e60b1b;
  wire al_e0e9a4f3;
  wire al_dbf8fa9d;
  wire al_f5f324f;
  wire al_6766b849;
  wire al_143e4872;
  wire al_a477b479;
  wire al_8bc3354;
  wire al_1e6bd6a1;
  wire al_e69868df;
  wire al_ae74b6ce;
  wire al_9290634f;
  wire al_7af9dc;
  wire al_8084b00c;
  wire al_b760f405;
  wire al_65d1cfc2;
  wire al_117e7922;
  wire al_633d0b30;
  wire al_b3570833;
  wire al_b9b8f3e1;
  wire al_37f2f859;
  wire al_691ab75e;
  wire al_78df4457;
  wire al_ea3d8437;
  wire al_d03ec855;
  wire al_d1805774;
  wire al_b2501f7c;
  wire al_2e361070;
  wire al_9b14b36d;
  wire al_e0fb24bc;
  wire al_2434069f;
  wire al_f06b68e;
  wire al_eed0f9b1;
  wire al_3fdcd506;
  wire al_8b101552;
  wire al_6d93b728;
  wire al_fef237c0;
  wire al_1a734e00;
  wire al_450062f6;
  wire al_96c7325f;
  wire al_34dcc703;
  wire al_8581252c;
  wire al_47ef5621;
  wire al_5595f015;
  wire al_7cd1dfe0;
  wire al_3baab685;
  wire al_bfe04e37;
  wire al_ff7baa95;
  wire al_4beff26f;
  wire al_215503f7;
  wire al_6ebcb190;
  wire al_e3b23b3d;
  wire al_27782d3b;
  wire al_96a09b29;
  wire al_f5c79977;
  wire al_d0973a8a;
  wire al_53ed7af5;
  wire al_f5a1ca8f;
  wire al_c40e7d13;
  wire al_b434c7b1;
  wire al_8d68d680;
  wire al_af211502;
  wire al_7b9dbd92;
  wire al_ce16dbbf;
  wire al_95f16875;
  wire al_81bff2a0;
  wire al_b661fbd8;
  wire al_d0b214a9;
  wire al_9fb02266;
  wire al_c2f2105d;
  wire al_df257acd;
  wire al_ceac5249;
  wire al_a09d4af8;
  wire al_8b2f2894;
  wire al_7ae76686;
  wire al_4d2bf11f;
  wire al_cedf3c10;
  wire al_4e77bfa;
  wire al_5efe66e3;
  wire al_693c6c75;
  wire al_822e59ab;
  wire al_5db6e161;
  wire al_34b35b3f;
  wire al_5010b887;
  wire al_7d8a00ee;
  wire al_9bd13530;
  wire al_a0c66e60;
  wire al_aab46c70;
  wire al_7b742de5;
  wire al_5b895c4d;
  wire al_8526f7d0;
  wire al_3dd7b884;
  wire al_9c8e7269;
  wire al_216fbee;
  wire al_fdd42739;
  wire al_ed1e8e02;
  wire al_8208c979;
  wire al_2842b1a1;
  wire al_594d587;
  wire al_f57392c;
  wire al_9dc8cf16;
  wire al_23f7cf96;
  wire al_6007eb01;
  wire al_e9dcbf51;
  wire al_af282b4e;
  wire al_f13375bf;
  wire al_79e6f53f;
  wire al_262f4fd9;
  wire al_91a1715;
  wire al_466678a0;
  wire al_b3412438;
  wire al_905abb5d;
  wire al_30d2d597;
  wire al_b4ebcfb5;
  wire al_9398f98d;
  wire al_2e77c07b;
  wire al_56c765b9;
  wire al_abeeae47;
  wire al_59c21146;
  wire al_e154cc8;
  wire al_c2370696;
  wire al_c0c45a44;
  wire al_32d5e65b;
  wire al_627e2733;
  wire al_4caf87a4;
  wire al_93eba83e;
  wire al_f4b95543;
  wire al_431d20ff;
  wire al_12da8cbc;
  wire al_a05b5ad4;
  wire al_5072fc21;
  wire al_e6b19e19;
  wire al_baadae4d;
  wire al_c4be0e1d;
  wire al_5dc8be80;
  wire al_547ff558;
  wire al_ecd1dd20;
  wire al_a4a9db62;
  wire al_2150e0ab;
  wire al_98763df0;
  wire al_a2aa2d49;
  wire al_e749a18b;
  wire al_65250a4c;
  wire al_71dba21f;
  wire al_5ba1798e;
  wire al_fa3cfc2c;
  wire al_eebdc4f4;
  wire al_88900ac6;
  wire al_f1ea9238;
  wire al_cb718520;
  wire al_47b988e0;
  wire al_919eb56e;
  wire al_35e6fce8;
  wire al_6a0855b2;
  wire al_607eee13;
  wire al_9f13bda9;
  wire al_7d943beb;
  wire al_6d747586;
  wire al_d6a2647c;
  wire al_8cb59e89;
  wire al_63e85dd3;
  wire al_2d304c84;
  wire al_59db63b2;
  wire al_ef9e6ec2;
  wire al_ee134d8c;
  wire al_931bfadf;
  wire al_f57240df;
  wire al_d1cf7fc7;
  wire al_f80ea3fa;
  wire al_6cebde96;
  wire al_4e2c20db;
  wire al_5334aacc;
  wire al_c6f75c3f;
  wire al_d26c1ceb;
  wire al_22bff0ea;
  wire al_38e51a5b;
  wire al_6b77e7f1;
  wire al_93915853;
  wire al_6abbbc54;
  wire al_aa70c10f;
  wire al_41b2a88c;
  wire al_dde17c7f;
  wire al_6df879f;
  wire al_ca3af73f;
  wire al_b8b96eac;
  wire al_d7300a25;
  wire al_9c595c5;
  wire al_b47bbe21;
  wire al_e295dc49;
  wire al_85e166c5;
  wire al_689afff7;
  wire al_36c0ab0e;
  wire al_9cf8f60d;
  wire al_a8352957;
  wire al_be007839;
  wire al_66995ad4;
  wire al_4dcb599e;
  wire al_155419a5;
  wire al_49b8db26;
  wire al_8468641;
  wire al_9f4fbb79;
  wire al_732042af;
  wire al_cd055708;
  wire al_2e4b86ef;
  wire al_b84db2a6;
  wire al_526f98e2;
  wire al_e6e3fffa;
  wire al_5b27964b;
  wire al_9459711;
  wire al_1fb17bb2;
  wire al_35fbae96;
  wire al_453ca3a4;
  wire al_e907e498;
  wire al_e1852c9f;
  wire al_3432ca06;
  wire al_41ebf214;
  wire al_57ac52e7;
  wire al_2b438376;
  wire al_ca3e9bc8;
  wire al_464b5ec;
  wire al_a0e81a0c;
  wire al_6e619896;
  wire al_f3664844;
  wire al_eb180f53;
  wire al_ad51aadd;
  wire al_aa6720b4;
  wire al_82c92bf1;
  wire al_51ccac31;
  wire al_a50d3ef5;
  wire al_b9439b67;
  wire al_24f0c9b4;
  wire al_8e479b1b;
  wire al_6aa12cb6;
  wire al_1d3f4f78;
  wire al_63e4776;
  wire al_fb5dab05;
  wire al_2e3e139;
  wire al_92d8d26e;
  wire al_94cd12cf;
  wire al_31ed294d;
  wire al_58d02051;
  wire al_1024d4fd;
  wire al_c1da9790;
  wire al_6cad4dc9;
  wire al_2abe7dd5;
  wire al_441d631;
  wire al_f3239c7d;
  wire al_b87907a9;
  wire al_90f0f7d8;
  wire al_a4b7f674;
  wire al_7076449e;
  wire al_8e44a4d6;
  wire al_4ff3fb03;
  wire al_724c9346;
  wire al_654ec6c7;
  wire al_db43acf6;
  wire al_1881b524;
  wire al_ee4e9a87;
  wire al_ea6aa5ed;
  wire al_d4f16200;
  wire al_ee99ca7f;
  wire al_b8f391da;
  wire al_98d4708b;
  wire al_e355574b;
  wire al_750642c9;
  wire al_ff2d726;
  wire al_53853e4b;
  wire al_89b35cc7;
  wire al_375b5a4d;
  wire al_12dcd287;
  wire al_ff1931b3;
  wire al_4bd1c0eb;
  wire al_ac55c9d9;
  wire al_869b4e37;
  wire al_ca5ea173;
  wire al_76985513;
  wire al_8b8db5a8;
  wire al_8d3dc6f8;
  wire al_af8cdc32;
  wire al_50432123;
  wire al_2637e6b1;
  wire al_d2ba203e;
  wire al_72aa54c;
  wire al_5c60fab;
  wire al_aa0aca8a;
  wire al_26b3b41e;
  wire al_27f44dd8;
  wire al_8b60a1f7;

  AL_DFF_X al_468ea82d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_51794c84),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3da4ff6f[0]));
  AL_DFF_X al_f05d54ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[46]));
  AL_DFF_X al_1b02ef40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[47]));
  AL_DFF_X al_aaf901a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[48]));
  AL_DFF_X al_2c28460a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[49]));
  AL_DFF_X al_8f61afcc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[50]));
  AL_DFF_X al_72ebfd98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[51]));
  AL_DFF_X al_96b47a47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[52]));
  AL_DFF_X al_9e968c91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[53]));
  AL_DFF_X al_6f9571f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[54]));
  AL_DFF_X al_9328869 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[55]));
  AL_DFF_X al_9501021e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[56]));
  AL_DFF_X al_b598af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[57]));
  AL_DFF_X al_c0f6a9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[58]));
  AL_DFF_X al_e4349418 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[59]));
  AL_DFF_X al_e70d611d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[60]));
  AL_DFF_X al_6ad4b247 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[61]));
  AL_DFF_X al_2095fdca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[62]));
  AL_DFF_X al_fef08054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[63]));
  AL_DFF_X al_5e257bd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[64]));
  AL_DFF_X al_31366301 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[65]));
  AL_DFF_X al_11f9ca66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[66]));
  AL_DFF_X al_e75a1427 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[67]));
  AL_DFF_X al_291aeb7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[68]));
  AL_DFF_X al_be427733 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[69]));
  AL_DFF_X al_4394dead (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[70]));
  AL_DFF_X al_b9260c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[71]));
  AL_DFF_X al_b5e3e14d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[72]));
  AL_DFF_X al_370111e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[73]));
  AL_DFF_X al_38252f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[74]));
  AL_DFF_X al_6e209dc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[75]));
  AL_DFF_X al_fe119f0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[76]));
  AL_DFF_X al_cbc577f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d1d5c0[78]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3bd314e4[77]));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(~E*D))"),
    .INIT(32'h80800080))
    al_7329fe53 (
    .a(al_56e18a80),
    .b(al_e0cc30a4),
    .c(al_e8aefc81),
    .d(al_9d1d5c0[47]),
    .e(al_a5806bc7[47]),
    .o(al_689ce8c2));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_fceac18b (
    .a(al_9d1d5c0[72]),
    .b(al_9d1d5c0[73]),
    .c(al_9d1d5c0[74]),
    .d(al_9d1d5c0[75]),
    .e(al_9d1d5c0[76]),
    .f(al_9d1d5c0[77]),
    .o(al_147773d6));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_7d20f6bd (
    .a(al_9d1d5c0[60]),
    .b(al_9d1d5c0[61]),
    .c(al_9d1d5c0[62]),
    .d(al_9d1d5c0[63]),
    .e(al_9d1d5c0[64]),
    .f(al_9d1d5c0[65]),
    .o(al_4a4b505));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_83ecb74b (
    .a(al_1e3141cc),
    .b(al_4a4b505),
    .c(al_9d1d5c0[48]),
    .d(al_9d1d5c0[49]),
    .e(al_9d1d5c0[50]),
    .f(al_9d1d5c0[51]),
    .o(al_e8aefc81));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*C*B*A))"),
    .INIT(32'h7fff0000))
    al_13708e22 (
    .a(al_56e18a80),
    .b(al_e0cc30a4),
    .c(al_e8aefc81),
    .d(al_9d1d5c0[47]),
    .e(al_a5806bc7[47]),
    .o(al_d3fd7d5a[47]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_e908180a (
    .a(al_147773d6),
    .b(al_9d1d5c0[78]),
    .o(al_56e18a80));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_71798e22 (
    .a(al_9d1d5c0[54]),
    .b(al_9d1d5c0[55]),
    .c(al_9d1d5c0[56]),
    .d(al_9d1d5c0[57]),
    .e(al_9d1d5c0[58]),
    .f(al_9d1d5c0[59]),
    .o(al_1435a49e));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_682c8b1 (
    .a(al_1435a49e),
    .b(al_9d1d5c0[52]),
    .c(al_9d1d5c0[53]),
    .o(al_e0cc30a4));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_9ac9a737 (
    .a(al_9d1d5c0[66]),
    .b(al_9d1d5c0[67]),
    .c(al_9d1d5c0[68]),
    .d(al_9d1d5c0[69]),
    .e(al_9d1d5c0[70]),
    .f(al_9d1d5c0[71]),
    .o(al_1e3141cc));
  AL_DFF_X al_4d678d84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[0]));
  AL_DFF_X al_2a67f561 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[9]));
  AL_DFF_X al_9f7da054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[10]));
  AL_DFF_X al_578a5e4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[11]));
  AL_DFF_X al_6fdef335 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[12]));
  AL_DFF_X al_b5e39760 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[13]));
  AL_DFF_X al_10b76c47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[14]));
  AL_DFF_X al_568b8612 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[15]));
  AL_DFF_X al_f5cde503 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[16]));
  AL_DFF_X al_15d0ac29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[17]));
  AL_DFF_X al_4884095a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[18]));
  AL_DFF_X al_fb3db78a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[1]));
  AL_DFF_X al_8c187e33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[19]));
  AL_DFF_X al_680065bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[20]));
  AL_DFF_X al_1cc571b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[21]));
  AL_DFF_X al_71a25c65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[22]));
  AL_DFF_X al_dbe49e61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[23]));
  AL_DFF_X al_720eed44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[24]));
  AL_DFF_X al_c16c18e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[25]));
  AL_DFF_X al_df4e0abc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[26]));
  AL_DFF_X al_2d55d85b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[27]));
  AL_DFF_X al_2ad4ec43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[28]));
  AL_DFF_X al_97cbd42f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[2]));
  AL_DFF_X al_aef212ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[29]));
  AL_DFF_X al_1d1de29f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[30]));
  AL_DFF_X al_4af6d0fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[31]));
  AL_DFF_X al_25baf6dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[32]));
  AL_DFF_X al_38a1541d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[33]));
  AL_DFF_X al_e041ede0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[34]));
  AL_DFF_X al_49ddd5e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[35]));
  AL_DFF_X al_809b1ccb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[36]));
  AL_DFF_X al_e3abfc0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[37]));
  AL_DFF_X al_902b36a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[38]));
  AL_DFF_X al_bec6e92d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[3]));
  AL_DFF_X al_fc0a19be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[39]));
  AL_DFF_X al_d7aa4532 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[40]));
  AL_DFF_X al_b0e53702 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[41]));
  AL_DFF_X al_989def08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[42]));
  AL_DFF_X al_955ed71d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[43]));
  AL_DFF_X al_c00141d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[44]));
  AL_DFF_X al_346077 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[45]));
  AL_DFF_X al_946c141 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[46]));
  AL_DFF_X al_afed33a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3fd7d5a[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[47]));
  AL_DFF_X al_cb6cd8b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[4]));
  AL_DFF_X al_a6193522 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[5]));
  AL_DFF_X al_c4c2575d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[6]));
  AL_DFF_X al_14cd5258 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[7]));
  AL_DFF_X al_b5245bc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5806bc7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_83a08f3f[8]));
  AL_DFF_X al_73ac1b5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_689ce8c2),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_33c3313d[0]));
  AL_DFF_X al_6152a3ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4b6a4daa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_adb04807[0]));
  AL_DFF_X al_5f79a6d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[36]));
  AL_DFF_X al_78e2057d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[37]));
  AL_DFF_X al_272e98b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[38]));
  AL_DFF_X al_965ccab7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[39]));
  AL_DFF_X al_a6526f53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[40]));
  AL_DFF_X al_81dd4528 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[41]));
  AL_DFF_X al_3b902de2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[42]));
  AL_DFF_X al_d1b64535 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[43]));
  AL_DFF_X al_a4b78cc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[44]));
  AL_DFF_X al_d94db645 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[45]));
  AL_DFF_X al_f2abe165 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[46]));
  AL_DFF_X al_49ab6140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[47]));
  AL_DFF_X al_641f795c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[48]));
  AL_DFF_X al_3e38d366 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[49]));
  AL_DFF_X al_df8c9b79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[50]));
  AL_DFF_X al_107d1a0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[51]));
  AL_DFF_X al_b8e7d9cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[52]));
  AL_DFF_X al_e7c7c6d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[53]));
  AL_DFF_X al_3b2cedfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[54]));
  AL_DFF_X al_d3114476 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[55]));
  AL_DFF_X al_e095f19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[56]));
  AL_DFF_X al_d93cfbf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[57]));
  AL_DFF_X al_29a0c2a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[58]));
  AL_DFF_X al_b7f5fe18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[59]));
  AL_DFF_X al_d4a93acc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[60]));
  AL_DFF_X al_3fcb85a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[61]));
  AL_DFF_X al_7d0919e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[62]));
  AL_DFF_X al_331effc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[63]));
  AL_DFF_X al_e8830353 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[64]));
  AL_DFF_X al_d57cd3c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[65]));
  AL_DFF_X al_2d702a8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[66]));
  AL_DFF_X al_d71f4ecf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6f9059d1[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_177a13cd[67]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_127078a8 (
    .a(1'b0),
    .o({al_b32218f4,open_n2}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ebc9378f (
    .a(al_f2b51288[37]),
    .b(al_6f9059d1[37]),
    .c(al_b32218f4),
    .o({al_aa787729,al_6a5d599[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17b8d69c (
    .a(al_f2b51288[38]),
    .b(al_6f9059d1[38]),
    .c(al_aa787729),
    .o({al_c9b85978,al_6a5d599[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b5f4650b (
    .a(al_f2b51288[39]),
    .b(al_6f9059d1[39]),
    .c(al_c9b85978),
    .o({al_1472bf2f,al_6a5d599[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_21c1dfd7 (
    .a(al_f2b51288[40]),
    .b(al_6f9059d1[40]),
    .c(al_1472bf2f),
    .o({al_787b0a64,al_6a5d599[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_350cb68c (
    .a(al_f2b51288[41]),
    .b(al_6f9059d1[41]),
    .c(al_787b0a64),
    .o({al_c3020830,al_6a5d599[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4d1e8f6c (
    .a(al_f2b51288[42]),
    .b(al_6f9059d1[42]),
    .c(al_c3020830),
    .o({al_fa8bcfd,al_6a5d599[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_859c521c (
    .a(al_f2b51288[43]),
    .b(al_6f9059d1[43]),
    .c(al_fa8bcfd),
    .o({al_258d6ce0,al_6a5d599[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17a6d7fa (
    .a(al_f2b51288[44]),
    .b(al_6f9059d1[44]),
    .c(al_258d6ce0),
    .o({al_dc10836c,al_6a5d599[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dc4c0a98 (
    .a(al_f2b51288[45]),
    .b(al_6f9059d1[45]),
    .c(al_dc10836c),
    .o({al_4de5b5ba,al_6a5d599[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c1b88eb9 (
    .a(al_f2b51288[46]),
    .b(al_6f9059d1[46]),
    .c(al_4de5b5ba),
    .o({al_1a08a0b7,al_6a5d599[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_13bce3bb (
    .a(al_f2b51288[47]),
    .b(al_6f9059d1[47]),
    .c(al_1a08a0b7),
    .o({al_fe80d5e5,al_6a5d599[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a8c0e3a7 (
    .c(al_fe80d5e5),
    .o({open_n5,al_6a5d599[11]}));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_a4f8cdb5 (
    .a(al_95c9121c),
    .b(al_6a5d599[0]),
    .c(al_f2b51288[37]),
    .o(al_5d497694[37]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_99d58474 (
    .a(al_95c9121c),
    .b(al_6a5d599[1]),
    .c(al_f2b51288[38]),
    .o(al_5d497694[38]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_5c366e3b (
    .a(al_6f9059d1[63]),
    .b(al_6f9059d1[64]),
    .c(al_6f9059d1[65]),
    .d(al_6f9059d1[66]),
    .e(al_6f9059d1[67]),
    .f(al_6f9059d1[68]),
    .o(al_56ca40b1));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_d06dcdd0 (
    .a(al_95c9121c),
    .b(al_6a5d599[2]),
    .c(al_f2b51288[39]),
    .o(al_5d497694[39]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_ca76153c (
    .a(al_6f9059d1[57]),
    .b(al_6f9059d1[58]),
    .c(al_6f9059d1[59]),
    .d(al_6f9059d1[60]),
    .e(al_6f9059d1[61]),
    .f(al_6f9059d1[62]),
    .o(al_2f2f061f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_627cd07 (
    .a(al_6f9059d1[51]),
    .b(al_6f9059d1[52]),
    .c(al_6f9059d1[53]),
    .d(al_6f9059d1[54]),
    .e(al_6f9059d1[55]),
    .f(al_6f9059d1[56]),
    .o(al_75e67c73));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_fdf9106b (
    .a(al_6a5d599[11]),
    .b(al_6f9059d1[48]),
    .c(al_6f9059d1[49]),
    .d(al_6f9059d1[50]),
    .o(al_93654000));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_517c054e (
    .a(al_56ca40b1),
    .b(al_2f2f061f),
    .c(al_75e67c73),
    .d(al_93654000),
    .o(al_95c9121c));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_43e58f39 (
    .a(al_95c9121c),
    .b(al_6a5d599[3]),
    .c(al_f2b51288[40]),
    .o(al_5d497694[40]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_4debe22a (
    .a(al_95c9121c),
    .b(al_6a5d599[4]),
    .c(al_f2b51288[41]),
    .o(al_5d497694[41]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_3de3f8d6 (
    .a(al_95c9121c),
    .b(al_6a5d599[5]),
    .c(al_f2b51288[42]),
    .o(al_5d497694[42]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_b16e2bba (
    .a(al_95c9121c),
    .b(al_6a5d599[6]),
    .c(al_f2b51288[43]),
    .o(al_5d497694[43]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_aa19c4f9 (
    .a(al_95c9121c),
    .b(al_6a5d599[7]),
    .c(al_f2b51288[44]),
    .o(al_5d497694[44]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_f0135bd9 (
    .a(al_95c9121c),
    .b(al_6a5d599[8]),
    .c(al_f2b51288[45]),
    .o(al_5d497694[45]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_5213dd26 (
    .a(al_95c9121c),
    .b(al_6a5d599[9]),
    .c(al_f2b51288[46]),
    .o(al_5d497694[46]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    al_9b9603e7 (
    .a(al_95c9121c),
    .b(al_6a5d599[10]),
    .c(al_f2b51288[47]),
    .o(al_5d497694[47]));
  AL_DFF_X al_8266a5e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[0]));
  AL_DFF_X al_1b49cda3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[9]));
  AL_DFF_X al_10a47e2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[10]));
  AL_DFF_X al_6b71d5f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[11]));
  AL_DFF_X al_ed7b70a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[12]));
  AL_DFF_X al_bd543057 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[13]));
  AL_DFF_X al_70345330 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[14]));
  AL_DFF_X al_b238e1c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[15]));
  AL_DFF_X al_73e64515 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[16]));
  AL_DFF_X al_7366212c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[17]));
  AL_DFF_X al_1b3562b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[18]));
  AL_DFF_X al_b1d8f7fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[1]));
  AL_DFF_X al_88ffef54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[19]));
  AL_DFF_X al_aa86b037 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[20]));
  AL_DFF_X al_c3eeb988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[21]));
  AL_DFF_X al_8f017b8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[22]));
  AL_DFF_X al_597ec2cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[23]));
  AL_DFF_X al_485a91ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[24]));
  AL_DFF_X al_6911f639 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[25]));
  AL_DFF_X al_555ae646 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[26]));
  AL_DFF_X al_134d895c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[27]));
  AL_DFF_X al_3628fbe2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[28]));
  AL_DFF_X al_18bbf4ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[2]));
  AL_DFF_X al_1325e582 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[29]));
  AL_DFF_X al_60a22d8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[30]));
  AL_DFF_X al_fcd51b04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[31]));
  AL_DFF_X al_65745020 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[32]));
  AL_DFF_X al_31fa29f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[33]));
  AL_DFF_X al_bbc287bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[34]));
  AL_DFF_X al_dfad6419 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[35]));
  AL_DFF_X al_4c57853c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[36]));
  AL_DFF_X al_dde22664 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[37]));
  AL_DFF_X al_b3992c97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[38]));
  AL_DFF_X al_20634034 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[3]));
  AL_DFF_X al_af2b2f29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[39]));
  AL_DFF_X al_9ba329d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[40]));
  AL_DFF_X al_c9b14a90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[41]));
  AL_DFF_X al_2eb435ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[42]));
  AL_DFF_X al_3212dcab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[43]));
  AL_DFF_X al_756cacb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[44]));
  AL_DFF_X al_173842c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[45]));
  AL_DFF_X al_d8fb36ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[46]));
  AL_DFF_X al_64e856b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d497694[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[47]));
  AL_DFF_X al_b8acecce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[4]));
  AL_DFF_X al_814952c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[5]));
  AL_DFF_X al_5f54b466 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[6]));
  AL_DFF_X al_e7634760 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[7]));
  AL_DFF_X al_aca4664 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2b51288[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6c6869d7[8]));
  AL_DFF_X al_2efb95f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_95c9121c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[0]));
  AL_DFF_X al_6bf49e2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[9]));
  AL_DFF_X al_5f3adf07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[10]));
  AL_DFF_X al_851e878d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[1]));
  AL_DFF_X al_964b1d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[2]));
  AL_DFF_X al_ea507f2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[3]));
  AL_DFF_X al_f19d90a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[4]));
  AL_DFF_X al_aafd4bab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[5]));
  AL_DFF_X al_62cf74c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[6]));
  AL_DFF_X al_5e2b635f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[7]));
  AL_DFF_X al_24495daf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fac191b8[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c9ed4b28[8]));
  AL_DFF_X al_d8b6cb2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_adb04807[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e1bd9dc[0]));
  AL_DFF_X al_6fae27d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[35]));
  AL_DFF_X al_1631ae61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[36]));
  AL_DFF_X al_beced3ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[37]));
  AL_DFF_X al_7b1c76ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[38]));
  AL_DFF_X al_5a79623b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[39]));
  AL_DFF_X al_a28b20f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[40]));
  AL_DFF_X al_a92bff3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[41]));
  AL_DFF_X al_cc5d3cff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[42]));
  AL_DFF_X al_d03fcb19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[43]));
  AL_DFF_X al_c1a312dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[44]));
  AL_DFF_X al_ec245c2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[45]));
  AL_DFF_X al_aaa171ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[46]));
  AL_DFF_X al_7ec2a1f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[47]));
  AL_DFF_X al_813959e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[48]));
  AL_DFF_X al_ea2dc1c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[49]));
  AL_DFF_X al_d102b7a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[50]));
  AL_DFF_X al_5f6e1db9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[51]));
  AL_DFF_X al_a8df7a3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[52]));
  AL_DFF_X al_da88ffc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[53]));
  AL_DFF_X al_7a8953eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[54]));
  AL_DFF_X al_ef619ade (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[55]));
  AL_DFF_X al_9178c76c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[56]));
  AL_DFF_X al_46f06370 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[57]));
  AL_DFF_X al_14b297f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[58]));
  AL_DFF_X al_fc7177c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[59]));
  AL_DFF_X al_a59e8436 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[60]));
  AL_DFF_X al_84a96949 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[61]));
  AL_DFF_X al_2f90f304 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[62]));
  AL_DFF_X al_e8fa0c7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[63]));
  AL_DFF_X al_54af62c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[64]));
  AL_DFF_X al_8c458ead (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[65]));
  AL_DFF_X al_a3f605dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_177a13cd[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a6f4a789[66]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_55467134 (
    .a(1'b0),
    .o({al_6a7cf4f6,open_n8}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a41f842a (
    .a(al_6c6869d7[36]),
    .b(al_177a13cd[36]),
    .c(al_6a7cf4f6),
    .o({al_7d43f9f9,al_2e720a5a[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_78b93eb8 (
    .a(al_6c6869d7[37]),
    .b(al_177a13cd[37]),
    .c(al_7d43f9f9),
    .o({al_c2244c00,al_2e720a5a[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bee03fed (
    .a(al_6c6869d7[38]),
    .b(al_177a13cd[38]),
    .c(al_c2244c00),
    .o({al_3690d0d4,al_2e720a5a[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c51efe30 (
    .a(al_6c6869d7[39]),
    .b(al_177a13cd[39]),
    .c(al_3690d0d4),
    .o({al_5b92a62d,al_2e720a5a[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d9d00c9f (
    .a(al_6c6869d7[40]),
    .b(al_177a13cd[40]),
    .c(al_5b92a62d),
    .o({al_59478e92,al_2e720a5a[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cba63229 (
    .a(al_6c6869d7[41]),
    .b(al_177a13cd[41]),
    .c(al_59478e92),
    .o({al_9ea91fcd,al_2e720a5a[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fbe9ae2d (
    .a(al_6c6869d7[42]),
    .b(al_177a13cd[42]),
    .c(al_9ea91fcd),
    .o({al_3d9987d2,al_2e720a5a[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2fad4cc3 (
    .a(al_6c6869d7[43]),
    .b(al_177a13cd[43]),
    .c(al_3d9987d2),
    .o({al_c5d02c43,al_2e720a5a[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f65f531c (
    .a(al_6c6869d7[44]),
    .b(al_177a13cd[44]),
    .c(al_c5d02c43),
    .o({al_8889fefd,al_2e720a5a[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a99991e (
    .a(al_6c6869d7[45]),
    .b(al_177a13cd[45]),
    .c(al_8889fefd),
    .o({al_28b0e45b,al_2e720a5a[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a15a1732 (
    .a(al_6c6869d7[46]),
    .b(al_177a13cd[46]),
    .c(al_28b0e45b),
    .o({al_1e2e550f,al_2e720a5a[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_74fb5b4d (
    .a(al_6c6869d7[47]),
    .b(al_177a13cd[47]),
    .c(al_1e2e550f),
    .o({al_3afa0b96,al_2e720a5a[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5a59f169 (
    .c(al_3afa0b96),
    .o({open_n11,al_2e720a5a[12]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d4cee76f (
    .a(al_82230b41),
    .b(al_6c6869d7[36]),
    .c(al_2e720a5a[0]),
    .o(al_c2901510[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9e1cf98d (
    .a(al_82230b41),
    .b(al_6c6869d7[37]),
    .c(al_2e720a5a[1]),
    .o(al_c2901510[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_71cbacc9 (
    .a(al_82230b41),
    .b(al_6c6869d7[38]),
    .c(al_2e720a5a[2]),
    .o(al_c2901510[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fb29e41d (
    .a(al_82230b41),
    .b(al_6c6869d7[39]),
    .c(al_2e720a5a[3]),
    .o(al_c2901510[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5a3eac91 (
    .a(al_82230b41),
    .b(al_6c6869d7[40]),
    .c(al_2e720a5a[4]),
    .o(al_c2901510[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_929b7aa4 (
    .a(al_82230b41),
    .b(al_6c6869d7[41]),
    .c(al_2e720a5a[5]),
    .o(al_c2901510[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4f047c65 (
    .a(al_82230b41),
    .b(al_6c6869d7[42]),
    .c(al_2e720a5a[6]),
    .o(al_c2901510[42]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_b1acb145 (
    .a(al_177a13cd[62]),
    .b(al_177a13cd[63]),
    .c(al_177a13cd[64]),
    .d(al_177a13cd[65]),
    .e(al_177a13cd[66]),
    .f(al_177a13cd[67]),
    .o(al_c029c247));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_589cfbd0 (
    .a(al_177a13cd[56]),
    .b(al_177a13cd[57]),
    .c(al_177a13cd[58]),
    .d(al_177a13cd[59]),
    .e(al_177a13cd[60]),
    .f(al_177a13cd[61]),
    .o(al_62aba81a));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_da6efe7b (
    .a(al_177a13cd[50]),
    .b(al_177a13cd[51]),
    .c(al_177a13cd[52]),
    .d(al_177a13cd[53]),
    .e(al_177a13cd[54]),
    .f(al_177a13cd[55]),
    .o(al_e889058f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*C*B*A)"),
    .INIT(64'h0000000000000080))
    al_122ea15f (
    .a(al_c029c247),
    .b(al_62aba81a),
    .c(al_e889058f),
    .d(al_177a13cd[48]),
    .e(al_177a13cd[49]),
    .f(al_2e720a5a[12]),
    .o(al_82230b41));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_626afeaf (
    .a(al_82230b41),
    .b(al_6c6869d7[43]),
    .c(al_2e720a5a[7]),
    .o(al_c2901510[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_63981119 (
    .a(al_82230b41),
    .b(al_6c6869d7[44]),
    .c(al_2e720a5a[8]),
    .o(al_c2901510[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d37187b8 (
    .a(al_82230b41),
    .b(al_6c6869d7[45]),
    .c(al_2e720a5a[9]),
    .o(al_c2901510[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ee126d43 (
    .a(al_82230b41),
    .b(al_6c6869d7[46]),
    .c(al_2e720a5a[10]),
    .o(al_c2901510[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1072140b (
    .a(al_82230b41),
    .b(al_6c6869d7[47]),
    .c(al_2e720a5a[11]),
    .o(al_c2901510[47]));
  AL_DFF_X al_ea63a970 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[0]));
  AL_DFF_X al_43388e59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[9]));
  AL_DFF_X al_f0d0ab77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[10]));
  AL_DFF_X al_9bdfd9db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[11]));
  AL_DFF_X al_8f6a70ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[12]));
  AL_DFF_X al_2d8c2d96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[13]));
  AL_DFF_X al_5c9c2c2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[14]));
  AL_DFF_X al_2d0decd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[15]));
  AL_DFF_X al_bcc45cd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[16]));
  AL_DFF_X al_eb02f765 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[17]));
  AL_DFF_X al_7bba172f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[18]));
  AL_DFF_X al_a223d7e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[1]));
  AL_DFF_X al_e5120449 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[19]));
  AL_DFF_X al_733c7bc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[20]));
  AL_DFF_X al_104259ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[21]));
  AL_DFF_X al_e0aea401 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[22]));
  AL_DFF_X al_7937606c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[23]));
  AL_DFF_X al_68b9d908 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[24]));
  AL_DFF_X al_ac54bd57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[25]));
  AL_DFF_X al_aca56c9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[26]));
  AL_DFF_X al_c4ed4ad9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[27]));
  AL_DFF_X al_66e89e91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[28]));
  AL_DFF_X al_390fbb5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[2]));
  AL_DFF_X al_7caa768a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[29]));
  AL_DFF_X al_5125691d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[30]));
  AL_DFF_X al_eb8690c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[31]));
  AL_DFF_X al_46d7739c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[32]));
  AL_DFF_X al_25c7ce1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[33]));
  AL_DFF_X al_23b41e78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[34]));
  AL_DFF_X al_cd66331a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[35]));
  AL_DFF_X al_71b4aafc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[36]));
  AL_DFF_X al_3e2be93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[37]));
  AL_DFF_X al_83c15d4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[38]));
  AL_DFF_X al_b624ce08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[3]));
  AL_DFF_X al_a079bc1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[39]));
  AL_DFF_X al_745002f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[40]));
  AL_DFF_X al_d6f15e9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[41]));
  AL_DFF_X al_af49a0b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[42]));
  AL_DFF_X al_b6b4fe2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[43]));
  AL_DFF_X al_f2743a70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[44]));
  AL_DFF_X al_2702263e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[45]));
  AL_DFF_X al_8a24188e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[46]));
  AL_DFF_X al_7039c2c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2901510[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[47]));
  AL_DFF_X al_b781f50d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[4]));
  AL_DFF_X al_343354b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[5]));
  AL_DFF_X al_d67df7df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[6]));
  AL_DFF_X al_4673131b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[7]));
  AL_DFF_X al_8ed4ed5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6c6869d7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d2e70f[8]));
  AL_DFF_X al_44537c05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82230b41),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[0]));
  AL_DFF_X al_4a95948c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[9]));
  AL_DFF_X al_884a8047 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[10]));
  AL_DFF_X al_6e606aef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[11]));
  AL_DFF_X al_82795640 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[1]));
  AL_DFF_X al_e31e4e2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[2]));
  AL_DFF_X al_88948916 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[3]));
  AL_DFF_X al_5894b362 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[4]));
  AL_DFF_X al_17145289 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[5]));
  AL_DFF_X al_d1c657d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[6]));
  AL_DFF_X al_136c7b82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[7]));
  AL_DFF_X al_b1b61de1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9ed4b28[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8fc8d46f[8]));
  AL_DFF_X al_9f488172 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e1bd9dc[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c6d10c98[0]));
  AL_DFF_X al_29fe0a73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[34]));
  AL_DFF_X al_23b2d88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[35]));
  AL_DFF_X al_5f542e81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[36]));
  AL_DFF_X al_a3abefef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[37]));
  AL_DFF_X al_8bd7ba75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[38]));
  AL_DFF_X al_2f43db1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[39]));
  AL_DFF_X al_f686383e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[40]));
  AL_DFF_X al_9058fff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[41]));
  AL_DFF_X al_3f69a20d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[42]));
  AL_DFF_X al_125abcc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[43]));
  AL_DFF_X al_3ab3918b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[44]));
  AL_DFF_X al_77591c8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[45]));
  AL_DFF_X al_72e69014 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[46]));
  AL_DFF_X al_e0f254bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[47]));
  AL_DFF_X al_74b92b74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[48]));
  AL_DFF_X al_b05cc67f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[49]));
  AL_DFF_X al_c837ff22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[50]));
  AL_DFF_X al_96e396cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[51]));
  AL_DFF_X al_a9562b1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[52]));
  AL_DFF_X al_147c51aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[53]));
  AL_DFF_X al_96b561fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[54]));
  AL_DFF_X al_af44bd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[55]));
  AL_DFF_X al_77bd78f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[56]));
  AL_DFF_X al_590f7421 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[57]));
  AL_DFF_X al_aba23386 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[58]));
  AL_DFF_X al_8049f251 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[59]));
  AL_DFF_X al_5454968 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[60]));
  AL_DFF_X al_aa92294a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[61]));
  AL_DFF_X al_67f0bbc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[62]));
  AL_DFF_X al_dbc46328 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[63]));
  AL_DFF_X al_9b53854a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[64]));
  AL_DFF_X al_bd912cdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a6f4a789[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_515b933[65]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_85f4c797 (
    .a(1'b0),
    .o({al_88df3967,open_n14}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c8a4deec (
    .a(al_13d2e70f[35]),
    .b(al_a6f4a789[35]),
    .c(al_88df3967),
    .o({al_2824b693,al_158480cc[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_daaacb7e (
    .a(al_13d2e70f[36]),
    .b(al_a6f4a789[36]),
    .c(al_2824b693),
    .o({al_6d794600,al_158480cc[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_adf58970 (
    .a(al_13d2e70f[37]),
    .b(al_a6f4a789[37]),
    .c(al_6d794600),
    .o({al_6e4bbf49,al_158480cc[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_28b00c77 (
    .a(al_13d2e70f[38]),
    .b(al_a6f4a789[38]),
    .c(al_6e4bbf49),
    .o({al_2ef9708,al_158480cc[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f1bbceff (
    .a(al_13d2e70f[39]),
    .b(al_a6f4a789[39]),
    .c(al_2ef9708),
    .o({al_f452a7c,al_158480cc[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_aa120909 (
    .a(al_13d2e70f[40]),
    .b(al_a6f4a789[40]),
    .c(al_f452a7c),
    .o({al_32e1725d,al_158480cc[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8d0014e1 (
    .a(al_13d2e70f[41]),
    .b(al_a6f4a789[41]),
    .c(al_32e1725d),
    .o({al_a83c9088,al_158480cc[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2d4215c2 (
    .a(al_13d2e70f[42]),
    .b(al_a6f4a789[42]),
    .c(al_a83c9088),
    .o({al_f9a74458,al_158480cc[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_702a4b45 (
    .a(al_13d2e70f[43]),
    .b(al_a6f4a789[43]),
    .c(al_f9a74458),
    .o({al_54803b10,al_158480cc[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_12836a8f (
    .a(al_13d2e70f[44]),
    .b(al_a6f4a789[44]),
    .c(al_54803b10),
    .o({al_7ba0f244,al_158480cc[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_23874c63 (
    .a(al_13d2e70f[45]),
    .b(al_a6f4a789[45]),
    .c(al_7ba0f244),
    .o({al_4e9b63c9,al_158480cc[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_db909ebf (
    .a(al_13d2e70f[46]),
    .b(al_a6f4a789[46]),
    .c(al_4e9b63c9),
    .o({al_dcea9b4,al_158480cc[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ce27dcc5 (
    .a(al_13d2e70f[47]),
    .b(al_a6f4a789[47]),
    .c(al_dcea9b4),
    .o({al_afad458d,al_158480cc[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9a685400 (
    .c(al_afad458d),
    .o({open_n17,al_158480cc[13]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_1d944862 (
    .a(al_a6f4a789[62]),
    .b(al_a6f4a789[63]),
    .c(al_a6f4a789[64]),
    .d(al_a6f4a789[65]),
    .e(al_a6f4a789[66]),
    .f(al_158480cc[13]),
    .o(al_90e336e1));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_d3306737 (
    .a(al_a6f4a789[56]),
    .b(al_a6f4a789[57]),
    .c(al_a6f4a789[58]),
    .d(al_a6f4a789[59]),
    .e(al_a6f4a789[60]),
    .f(al_a6f4a789[61]),
    .o(al_d41ac52e));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_22b5fef0 (
    .a(al_a6f4a789[50]),
    .b(al_a6f4a789[51]),
    .c(al_a6f4a789[52]),
    .d(al_a6f4a789[53]),
    .e(al_a6f4a789[54]),
    .f(al_a6f4a789[55]),
    .o(al_2bfcf033));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    al_d446af00 (
    .a(al_90e336e1),
    .b(al_d41ac52e),
    .c(al_2bfcf033),
    .d(al_a6f4a789[48]),
    .e(al_a6f4a789[49]),
    .o(al_bf8f4b75));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9fbc2c13 (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[35]),
    .c(al_158480cc[0]),
    .o(al_fb9cdc0e[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_664714d5 (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[36]),
    .c(al_158480cc[1]),
    .o(al_fb9cdc0e[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_873d04dd (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[37]),
    .c(al_158480cc[2]),
    .o(al_fb9cdc0e[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1c74cc33 (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[38]),
    .c(al_158480cc[3]),
    .o(al_fb9cdc0e[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8ec2ac01 (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[39]),
    .c(al_158480cc[4]),
    .o(al_fb9cdc0e[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_71e98eb4 (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[40]),
    .c(al_158480cc[5]),
    .o(al_fb9cdc0e[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ed210fe2 (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[41]),
    .c(al_158480cc[6]),
    .o(al_fb9cdc0e[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ed811ecb (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[42]),
    .c(al_158480cc[7]),
    .o(al_fb9cdc0e[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1e1fe231 (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[43]),
    .c(al_158480cc[8]),
    .o(al_fb9cdc0e[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_61efe8c (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[44]),
    .c(al_158480cc[9]),
    .o(al_fb9cdc0e[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2f17f8a9 (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[45]),
    .c(al_158480cc[10]),
    .o(al_fb9cdc0e[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2a789cf5 (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[46]),
    .c(al_158480cc[11]),
    .o(al_fb9cdc0e[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2110f6ae (
    .a(al_bf8f4b75),
    .b(al_13d2e70f[47]),
    .c(al_158480cc[12]),
    .o(al_fb9cdc0e[47]));
  AL_DFF_X al_f410e11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[0]));
  AL_DFF_X al_a016ed04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[9]));
  AL_DFF_X al_9e0ec8b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[10]));
  AL_DFF_X al_a565451c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[11]));
  AL_DFF_X al_be128d75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[12]));
  AL_DFF_X al_b2bf1119 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[13]));
  AL_DFF_X al_70174b36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[14]));
  AL_DFF_X al_94f45f23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[15]));
  AL_DFF_X al_328545 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[16]));
  AL_DFF_X al_d617d90d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[17]));
  AL_DFF_X al_d0cd4b9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[18]));
  AL_DFF_X al_26f7de1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[1]));
  AL_DFF_X al_7e7f3867 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[19]));
  AL_DFF_X al_df7c1c11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[20]));
  AL_DFF_X al_7db45bc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[21]));
  AL_DFF_X al_e2f7d4a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[22]));
  AL_DFF_X al_c8a2d143 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[23]));
  AL_DFF_X al_c02ced2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[24]));
  AL_DFF_X al_40f6285f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[25]));
  AL_DFF_X al_4071f2c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[26]));
  AL_DFF_X al_60ae7c64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[27]));
  AL_DFF_X al_85ff690c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[28]));
  AL_DFF_X al_8cd5ab0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[2]));
  AL_DFF_X al_f210341f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[29]));
  AL_DFF_X al_14c6601e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[30]));
  AL_DFF_X al_5196817f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[31]));
  AL_DFF_X al_12fcf706 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[32]));
  AL_DFF_X al_12a91d64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[33]));
  AL_DFF_X al_d926b261 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[34]));
  AL_DFF_X al_aeda6228 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[35]));
  AL_DFF_X al_cb015b59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[36]));
  AL_DFF_X al_6e92c339 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[37]));
  AL_DFF_X al_2b37ecde (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[38]));
  AL_DFF_X al_60029fa0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[3]));
  AL_DFF_X al_5c40e64e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[39]));
  AL_DFF_X al_d9c9a7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[40]));
  AL_DFF_X al_26f624dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[41]));
  AL_DFF_X al_ba9f6334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[42]));
  AL_DFF_X al_546ffbcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[43]));
  AL_DFF_X al_51ac833f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[44]));
  AL_DFF_X al_be5cc7b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[45]));
  AL_DFF_X al_f605efb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[46]));
  AL_DFF_X al_9bb9a4b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fb9cdc0e[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[47]));
  AL_DFF_X al_961aba1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[4]));
  AL_DFF_X al_27f54b2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[5]));
  AL_DFF_X al_8341a349 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[6]));
  AL_DFF_X al_b26f2647 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[7]));
  AL_DFF_X al_150a76b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d2e70f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7cada4c1[8]));
  AL_DFF_X al_d8eb92dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf8f4b75),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[0]));
  AL_DFF_X al_5c5f3a6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[9]));
  AL_DFF_X al_3a2f5421 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[10]));
  AL_DFF_X al_ea6471b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[11]));
  AL_DFF_X al_e3e71a5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[12]));
  AL_DFF_X al_91605568 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[1]));
  AL_DFF_X al_b0df883 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[2]));
  AL_DFF_X al_c25e4d28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[3]));
  AL_DFF_X al_e1b3426 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[4]));
  AL_DFF_X al_4c1f9ee5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[5]));
  AL_DFF_X al_22fe182f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[6]));
  AL_DFF_X al_2d229a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[7]));
  AL_DFF_X al_ac6b7e21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8fc8d46f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a63aa325[8]));
  AL_DFF_X al_21fc362f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c6d10c98[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_599810dd[0]));
  AL_DFF_X al_906d7fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[33]));
  AL_DFF_X al_a9c8640f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[34]));
  AL_DFF_X al_ec8cccaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[35]));
  AL_DFF_X al_95ac8f52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[36]));
  AL_DFF_X al_2e31fd1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[37]));
  AL_DFF_X al_b732c32d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[38]));
  AL_DFF_X al_f7a32431 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[39]));
  AL_DFF_X al_940491e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[40]));
  AL_DFF_X al_f551a605 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[41]));
  AL_DFF_X al_c9fc87ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[42]));
  AL_DFF_X al_68b50ac2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[43]));
  AL_DFF_X al_adbbef35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[44]));
  AL_DFF_X al_fe4ea5c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[45]));
  AL_DFF_X al_7138fafc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[46]));
  AL_DFF_X al_7f5221a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[47]));
  AL_DFF_X al_ae769e28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[48]));
  AL_DFF_X al_6850c9e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[49]));
  AL_DFF_X al_199c51bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[50]));
  AL_DFF_X al_e637da26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[51]));
  AL_DFF_X al_11e2235f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[52]));
  AL_DFF_X al_7c0ac2ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[53]));
  AL_DFF_X al_34f9f44b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[54]));
  AL_DFF_X al_d31a149a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[55]));
  AL_DFF_X al_f6cb0e34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[56]));
  AL_DFF_X al_56e5ee97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[57]));
  AL_DFF_X al_c887c678 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[58]));
  AL_DFF_X al_618bed49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[59]));
  AL_DFF_X al_3036169f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[60]));
  AL_DFF_X al_e180ca30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[61]));
  AL_DFF_X al_8eae9904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[62]));
  AL_DFF_X al_497e503f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[63]));
  AL_DFF_X al_9e385462 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_515b933[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_82ca84f8[64]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_40b88134 (
    .a(1'b0),
    .o({al_98398e18,open_n20}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a08bfd6 (
    .a(al_7cada4c1[34]),
    .b(al_515b933[34]),
    .c(al_98398e18),
    .o({al_463946df,al_4f616992[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6ba50150 (
    .a(al_7cada4c1[35]),
    .b(al_515b933[35]),
    .c(al_463946df),
    .o({al_967a5f00,al_4f616992[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3ccd5e9d (
    .a(al_7cada4c1[36]),
    .b(al_515b933[36]),
    .c(al_967a5f00),
    .o({al_110841cf,al_4f616992[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c1f0932c (
    .a(al_7cada4c1[37]),
    .b(al_515b933[37]),
    .c(al_110841cf),
    .o({al_9bebb94b,al_4f616992[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_baed19e8 (
    .a(al_7cada4c1[38]),
    .b(al_515b933[38]),
    .c(al_9bebb94b),
    .o({al_e2402cc4,al_4f616992[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b24d13e (
    .a(al_7cada4c1[39]),
    .b(al_515b933[39]),
    .c(al_e2402cc4),
    .o({al_49617358,al_4f616992[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd1e82de (
    .a(al_7cada4c1[40]),
    .b(al_515b933[40]),
    .c(al_49617358),
    .o({al_f9d08351,al_4f616992[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_890d5a7a (
    .a(al_7cada4c1[41]),
    .b(al_515b933[41]),
    .c(al_f9d08351),
    .o({al_57db75f0,al_4f616992[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_32ec2317 (
    .a(al_7cada4c1[42]),
    .b(al_515b933[42]),
    .c(al_57db75f0),
    .o({al_b261805d,al_4f616992[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3c7a0ff7 (
    .a(al_7cada4c1[43]),
    .b(al_515b933[43]),
    .c(al_b261805d),
    .o({al_d2377beb,al_4f616992[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b3f6820d (
    .a(al_7cada4c1[44]),
    .b(al_515b933[44]),
    .c(al_d2377beb),
    .o({al_f58e7482,al_4f616992[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_acf86999 (
    .a(al_7cada4c1[45]),
    .b(al_515b933[45]),
    .c(al_f58e7482),
    .o({al_2576177,al_4f616992[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a205ee1b (
    .a(al_7cada4c1[46]),
    .b(al_515b933[46]),
    .c(al_2576177),
    .o({al_64c2879,al_4f616992[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_546ed19c (
    .a(al_7cada4c1[47]),
    .b(al_515b933[47]),
    .c(al_64c2879),
    .o({al_6b5869dc,al_4f616992[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_98b4f76e (
    .c(al_6b5869dc),
    .o({open_n23,al_4f616992[14]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f12ba9c9 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[34]),
    .c(al_4f616992[0]),
    .o(al_28d525d8[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_958f37e9 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[35]),
    .c(al_4f616992[1]),
    .o(al_28d525d8[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b6248a18 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[36]),
    .c(al_4f616992[2]),
    .o(al_28d525d8[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3b934cd6 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[37]),
    .c(al_4f616992[3]),
    .o(al_28d525d8[37]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_4aa4106a (
    .a(al_515b933[60]),
    .b(al_515b933[61]),
    .c(al_515b933[62]),
    .d(al_515b933[63]),
    .e(al_515b933[64]),
    .f(al_515b933[65]),
    .o(al_f6f2dce7));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_ba1c2eff (
    .a(al_515b933[54]),
    .b(al_515b933[55]),
    .c(al_515b933[56]),
    .d(al_515b933[57]),
    .e(al_515b933[58]),
    .f(al_515b933[59]),
    .o(al_9cb945d3));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_1acff3ad (
    .a(al_515b933[48]),
    .b(al_515b933[49]),
    .c(al_515b933[50]),
    .d(al_515b933[51]),
    .e(al_515b933[52]),
    .f(al_515b933[53]),
    .o(al_c0342edb));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    al_6f7290db (
    .a(al_f6f2dce7),
    .b(al_9cb945d3),
    .c(al_c0342edb),
    .d(al_4f616992[14]),
    .o(al_abf1ad7c));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bdaedd42 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[38]),
    .c(al_4f616992[4]),
    .o(al_28d525d8[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_53ecba48 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[39]),
    .c(al_4f616992[5]),
    .o(al_28d525d8[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_eb3dcbf9 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[40]),
    .c(al_4f616992[6]),
    .o(al_28d525d8[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8d2cef72 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[41]),
    .c(al_4f616992[7]),
    .o(al_28d525d8[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1ae69b25 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[42]),
    .c(al_4f616992[8]),
    .o(al_28d525d8[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1acd4b73 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[43]),
    .c(al_4f616992[9]),
    .o(al_28d525d8[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f9a01bd5 (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[44]),
    .c(al_4f616992[10]),
    .o(al_28d525d8[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_17eadcd (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[45]),
    .c(al_4f616992[11]),
    .o(al_28d525d8[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cb357c0a (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[46]),
    .c(al_4f616992[12]),
    .o(al_28d525d8[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4582695d (
    .a(al_abf1ad7c),
    .b(al_7cada4c1[47]),
    .c(al_4f616992[13]),
    .o(al_28d525d8[47]));
  AL_DFF_X al_4616e159 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[0]));
  AL_DFF_X al_a542753a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[9]));
  AL_DFF_X al_60b64b90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[10]));
  AL_DFF_X al_94ff0074 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[11]));
  AL_DFF_X al_85ccce21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[12]));
  AL_DFF_X al_77102143 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[13]));
  AL_DFF_X al_bd32c96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[14]));
  AL_DFF_X al_245ff2ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[15]));
  AL_DFF_X al_6a75c46b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[16]));
  AL_DFF_X al_d7ce5939 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[17]));
  AL_DFF_X al_6c81427f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[18]));
  AL_DFF_X al_3ef3c680 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[1]));
  AL_DFF_X al_1a007d79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[19]));
  AL_DFF_X al_cd53d009 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[20]));
  AL_DFF_X al_417c7631 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[21]));
  AL_DFF_X al_2f3aea2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[22]));
  AL_DFF_X al_b4eabc45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[23]));
  AL_DFF_X al_325e5d4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[24]));
  AL_DFF_X al_8867859 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[25]));
  AL_DFF_X al_abc19d95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[26]));
  AL_DFF_X al_2cac10a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[27]));
  AL_DFF_X al_e29ad501 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[28]));
  AL_DFF_X al_fa562aaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[2]));
  AL_DFF_X al_a3063878 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[29]));
  AL_DFF_X al_95ffb542 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[30]));
  AL_DFF_X al_8c0b4207 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[31]));
  AL_DFF_X al_cdfdd29f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[32]));
  AL_DFF_X al_b4158b58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[33]));
  AL_DFF_X al_51ddb167 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[34]));
  AL_DFF_X al_83f4ae25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[35]));
  AL_DFF_X al_563dbc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[36]));
  AL_DFF_X al_56462c21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[37]));
  AL_DFF_X al_ee3e9548 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[38]));
  AL_DFF_X al_e118f7e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[3]));
  AL_DFF_X al_9fe4df51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[39]));
  AL_DFF_X al_f0375411 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[40]));
  AL_DFF_X al_11539140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[41]));
  AL_DFF_X al_8a9464b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[42]));
  AL_DFF_X al_67ff20c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[43]));
  AL_DFF_X al_e63e27a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[44]));
  AL_DFF_X al_5534f5b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[45]));
  AL_DFF_X al_9bf1600e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[46]));
  AL_DFF_X al_906a0916 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28d525d8[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[47]));
  AL_DFF_X al_3a757f27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[4]));
  AL_DFF_X al_71333c79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[5]));
  AL_DFF_X al_8f286034 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[6]));
  AL_DFF_X al_d49ae2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[7]));
  AL_DFF_X al_9dc6dc07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7cada4c1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5fd65077[8]));
  AL_DFF_X al_1e00f4e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abf1ad7c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[0]));
  AL_DFF_X al_b19d14db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[9]));
  AL_DFF_X al_92b46a58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[10]));
  AL_DFF_X al_1414e8a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[11]));
  AL_DFF_X al_affc17d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[12]));
  AL_DFF_X al_f57ab4ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[13]));
  AL_DFF_X al_a1773baf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[1]));
  AL_DFF_X al_dca95400 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[2]));
  AL_DFF_X al_7a3e34db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[3]));
  AL_DFF_X al_c4eb0b5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[4]));
  AL_DFF_X al_f4ce6afd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[5]));
  AL_DFF_X al_dd903039 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[6]));
  AL_DFF_X al_264c5a01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[7]));
  AL_DFF_X al_5b03cda2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a63aa325[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1898703d[8]));
  AL_DFF_X al_72c023ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_599810dd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_903e8807[0]));
  AL_DFF_X al_b3ec2850 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[32]));
  AL_DFF_X al_11ff4e46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[33]));
  AL_DFF_X al_a47b60ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[34]));
  AL_DFF_X al_1b148ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[35]));
  AL_DFF_X al_f3950344 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[36]));
  AL_DFF_X al_fb4994a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[37]));
  AL_DFF_X al_c230e97f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[38]));
  AL_DFF_X al_f48ee826 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[39]));
  AL_DFF_X al_1222aa4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[40]));
  AL_DFF_X al_6c98c7b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[41]));
  AL_DFF_X al_fcc4e257 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[42]));
  AL_DFF_X al_9dba4e0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[43]));
  AL_DFF_X al_b41d851e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[44]));
  AL_DFF_X al_8268c6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[45]));
  AL_DFF_X al_811df023 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[46]));
  AL_DFF_X al_98dc8c2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[47]));
  AL_DFF_X al_59d4b838 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[48]));
  AL_DFF_X al_e8b65af8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[49]));
  AL_DFF_X al_36be974 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[50]));
  AL_DFF_X al_74671485 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[51]));
  AL_DFF_X al_e9be3d34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[52]));
  AL_DFF_X al_2940be41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[53]));
  AL_DFF_X al_173a904b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[54]));
  AL_DFF_X al_e85f0701 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[55]));
  AL_DFF_X al_af52f041 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[56]));
  AL_DFF_X al_e90a2976 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[57]));
  AL_DFF_X al_59bd816f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[58]));
  AL_DFF_X al_4314159b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[59]));
  AL_DFF_X al_9fb8dba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[60]));
  AL_DFF_X al_fd09475b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[61]));
  AL_DFF_X al_accc1aae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[62]));
  AL_DFF_X al_d5ccc4a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_82ca84f8[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_297c219f[63]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_ba436f15 (
    .a(1'b0),
    .o({al_3971206e,open_n26}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cfbdc8fd (
    .a(al_5fd65077[33]),
    .b(al_82ca84f8[33]),
    .c(al_3971206e),
    .o({al_36535fd3,al_e67d7d00[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4515da29 (
    .a(al_5fd65077[34]),
    .b(al_82ca84f8[34]),
    .c(al_36535fd3),
    .o({al_430e5cec,al_e67d7d00[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_26b8737f (
    .a(al_5fd65077[35]),
    .b(al_82ca84f8[35]),
    .c(al_430e5cec),
    .o({al_35bf8c77,al_e67d7d00[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_401e0891 (
    .a(al_5fd65077[36]),
    .b(al_82ca84f8[36]),
    .c(al_35bf8c77),
    .o({al_6a165344,al_e67d7d00[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e996900c (
    .a(al_5fd65077[37]),
    .b(al_82ca84f8[37]),
    .c(al_6a165344),
    .o({al_edeaa856,al_e67d7d00[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_acff63b3 (
    .a(al_5fd65077[38]),
    .b(al_82ca84f8[38]),
    .c(al_edeaa856),
    .o({al_f3dfd21a,al_e67d7d00[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cf124edc (
    .a(al_5fd65077[39]),
    .b(al_82ca84f8[39]),
    .c(al_f3dfd21a),
    .o({al_b398ed4f,al_e67d7d00[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ad07bdd3 (
    .a(al_5fd65077[40]),
    .b(al_82ca84f8[40]),
    .c(al_b398ed4f),
    .o({al_5c1aec80,al_e67d7d00[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_775fa47a (
    .a(al_5fd65077[41]),
    .b(al_82ca84f8[41]),
    .c(al_5c1aec80),
    .o({al_1c3eecd0,al_e67d7d00[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bb0989a0 (
    .a(al_5fd65077[42]),
    .b(al_82ca84f8[42]),
    .c(al_1c3eecd0),
    .o({al_62e1f39,al_e67d7d00[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_44d3ca53 (
    .a(al_5fd65077[43]),
    .b(al_82ca84f8[43]),
    .c(al_62e1f39),
    .o({al_ee6cfa1b,al_e67d7d00[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f5789861 (
    .a(al_5fd65077[44]),
    .b(al_82ca84f8[44]),
    .c(al_ee6cfa1b),
    .o({al_7e84b0e7,al_e67d7d00[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4b2995a (
    .a(al_5fd65077[45]),
    .b(al_82ca84f8[45]),
    .c(al_7e84b0e7),
    .o({al_36b609cf,al_e67d7d00[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2d8dd4ed (
    .a(al_5fd65077[46]),
    .b(al_82ca84f8[46]),
    .c(al_36b609cf),
    .o({al_e216e162,al_e67d7d00[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2aecc401 (
    .a(al_5fd65077[47]),
    .b(al_82ca84f8[47]),
    .c(al_e216e162),
    .o({al_436534ab,al_e67d7d00[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_23d99bf (
    .c(al_436534ab),
    .o({open_n29,al_e67d7d00[15]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_961a02b2 (
    .a(al_ca0bc000),
    .b(al_5fd65077[33]),
    .c(al_e67d7d00[0]),
    .o(al_8d341179[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a6579192 (
    .a(al_ca0bc000),
    .b(al_5fd65077[34]),
    .c(al_e67d7d00[1]),
    .o(al_8d341179[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bc0ce376 (
    .a(al_ca0bc000),
    .b(al_5fd65077[35]),
    .c(al_e67d7d00[2]),
    .o(al_8d341179[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_edd675aa (
    .a(al_ca0bc000),
    .b(al_5fd65077[36]),
    .c(al_e67d7d00[3]),
    .o(al_8d341179[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_55ea699b (
    .a(al_ca0bc000),
    .b(al_5fd65077[37]),
    .c(al_e67d7d00[4]),
    .o(al_8d341179[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4213e9f5 (
    .a(al_ca0bc000),
    .b(al_5fd65077[38]),
    .c(al_e67d7d00[5]),
    .o(al_8d341179[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ec8ecf78 (
    .a(al_ca0bc000),
    .b(al_5fd65077[39]),
    .c(al_e67d7d00[6]),
    .o(al_8d341179[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_caae3e48 (
    .a(al_ca0bc000),
    .b(al_5fd65077[40]),
    .c(al_e67d7d00[7]),
    .o(al_8d341179[40]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_9dbef731 (
    .a(al_82ca84f8[60]),
    .b(al_82ca84f8[61]),
    .c(al_82ca84f8[62]),
    .d(al_82ca84f8[63]),
    .e(al_82ca84f8[64]),
    .f(al_e67d7d00[15]),
    .o(al_1a52e2b9));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_173b557 (
    .a(al_82ca84f8[54]),
    .b(al_82ca84f8[55]),
    .c(al_82ca84f8[56]),
    .d(al_82ca84f8[57]),
    .e(al_82ca84f8[58]),
    .f(al_82ca84f8[59]),
    .o(al_1686893d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_4dd493bc (
    .a(al_82ca84f8[48]),
    .b(al_82ca84f8[49]),
    .c(al_82ca84f8[50]),
    .d(al_82ca84f8[51]),
    .e(al_82ca84f8[52]),
    .f(al_82ca84f8[53]),
    .o(al_8c362b8c));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_b19f050d (
    .a(al_1a52e2b9),
    .b(al_1686893d),
    .c(al_8c362b8c),
    .o(al_ca0bc000));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d4339822 (
    .a(al_ca0bc000),
    .b(al_5fd65077[41]),
    .c(al_e67d7d00[8]),
    .o(al_8d341179[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b1aeba08 (
    .a(al_ca0bc000),
    .b(al_5fd65077[42]),
    .c(al_e67d7d00[9]),
    .o(al_8d341179[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_20dd76b0 (
    .a(al_ca0bc000),
    .b(al_5fd65077[43]),
    .c(al_e67d7d00[10]),
    .o(al_8d341179[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_49476ccb (
    .a(al_ca0bc000),
    .b(al_5fd65077[44]),
    .c(al_e67d7d00[11]),
    .o(al_8d341179[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9a4b835b (
    .a(al_ca0bc000),
    .b(al_5fd65077[45]),
    .c(al_e67d7d00[12]),
    .o(al_8d341179[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c75b0d5c (
    .a(al_ca0bc000),
    .b(al_5fd65077[46]),
    .c(al_e67d7d00[13]),
    .o(al_8d341179[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fbad1629 (
    .a(al_ca0bc000),
    .b(al_5fd65077[47]),
    .c(al_e67d7d00[14]),
    .o(al_8d341179[47]));
  AL_DFF_X al_e39c3db5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[0]));
  AL_DFF_X al_f025b104 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[9]));
  AL_DFF_X al_963c81b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[10]));
  AL_DFF_X al_59d09113 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[11]));
  AL_DFF_X al_91ec7cd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[12]));
  AL_DFF_X al_cb41e6fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[13]));
  AL_DFF_X al_1a6b3679 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[14]));
  AL_DFF_X al_e648e6ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[15]));
  AL_DFF_X al_91205465 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[16]));
  AL_DFF_X al_75ac6d43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[17]));
  AL_DFF_X al_9d156c4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[18]));
  AL_DFF_X al_3ae2830 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[1]));
  AL_DFF_X al_b4c3e574 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[19]));
  AL_DFF_X al_5176e269 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[20]));
  AL_DFF_X al_9866966f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[21]));
  AL_DFF_X al_14bda149 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[22]));
  AL_DFF_X al_df5ca051 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[23]));
  AL_DFF_X al_85e668ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[24]));
  AL_DFF_X al_510a1d16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[25]));
  AL_DFF_X al_363ce036 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[26]));
  AL_DFF_X al_3f1a3433 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[27]));
  AL_DFF_X al_542b48e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[28]));
  AL_DFF_X al_2cee7aa2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[2]));
  AL_DFF_X al_99518a8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[29]));
  AL_DFF_X al_c5608779 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[30]));
  AL_DFF_X al_920d907e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[31]));
  AL_DFF_X al_a6249348 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[32]));
  AL_DFF_X al_116b259a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[33]));
  AL_DFF_X al_64f67cbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[34]));
  AL_DFF_X al_643bb5d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[35]));
  AL_DFF_X al_33a30fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[36]));
  AL_DFF_X al_682c89a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[37]));
  AL_DFF_X al_41f7b64b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[38]));
  AL_DFF_X al_a95f4295 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[3]));
  AL_DFF_X al_58b8d7f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[39]));
  AL_DFF_X al_6af01a3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[40]));
  AL_DFF_X al_e5f2f3d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[41]));
  AL_DFF_X al_65665f5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[42]));
  AL_DFF_X al_e51a91f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[43]));
  AL_DFF_X al_ec9f70f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[44]));
  AL_DFF_X al_cf2b6dbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[45]));
  AL_DFF_X al_d2bf7219 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[46]));
  AL_DFF_X al_58a302fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d341179[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[47]));
  AL_DFF_X al_a4c63a08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[4]));
  AL_DFF_X al_664bbff3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[5]));
  AL_DFF_X al_e092d1cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[6]));
  AL_DFF_X al_69d841a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[7]));
  AL_DFF_X al_bd9a3cfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5fd65077[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_174c5039[8]));
  AL_DFF_X al_bc3082cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ca0bc000),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[0]));
  AL_DFF_X al_517a5fb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[9]));
  AL_DFF_X al_ac709ec3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[10]));
  AL_DFF_X al_e64b0190 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[11]));
  AL_DFF_X al_fd4813f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[12]));
  AL_DFF_X al_46e114bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[13]));
  AL_DFF_X al_5fc29a39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[14]));
  AL_DFF_X al_8d947be7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[1]));
  AL_DFF_X al_9eb67271 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[2]));
  AL_DFF_X al_1808ee31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[3]));
  AL_DFF_X al_51f91994 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[4]));
  AL_DFF_X al_f5d4682f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[5]));
  AL_DFF_X al_4f892e5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[6]));
  AL_DFF_X al_790c5e6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[7]));
  AL_DFF_X al_f63cccb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1898703d[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ebfa785c[8]));
  AL_DFF_X al_a7134794 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_903e8807[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5ed5f44b[0]));
  AL_DFF_X al_35729cab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[31]));
  AL_DFF_X al_d8477bfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[32]));
  AL_DFF_X al_6b8fc532 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[33]));
  AL_DFF_X al_e30f50e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[34]));
  AL_DFF_X al_d749ac03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[35]));
  AL_DFF_X al_577090d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[36]));
  AL_DFF_X al_f2f0538b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[37]));
  AL_DFF_X al_1d78249 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[38]));
  AL_DFF_X al_3abe078b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[39]));
  AL_DFF_X al_722c2ab2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[40]));
  AL_DFF_X al_14f30929 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[41]));
  AL_DFF_X al_e85ffc3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[42]));
  AL_DFF_X al_ab41cdcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[43]));
  AL_DFF_X al_f3cee596 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[44]));
  AL_DFF_X al_45fd4996 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[45]));
  AL_DFF_X al_506666b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[46]));
  AL_DFF_X al_6b2aea0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[47]));
  AL_DFF_X al_d15409ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[48]));
  AL_DFF_X al_605d89f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[49]));
  AL_DFF_X al_ac0385bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[50]));
  AL_DFF_X al_a5e4ca0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[51]));
  AL_DFF_X al_73a80b63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[52]));
  AL_DFF_X al_6b8e72e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[53]));
  AL_DFF_X al_6fedd4db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[54]));
  AL_DFF_X al_2ec6a9ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[55]));
  AL_DFF_X al_fc6653ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[56]));
  AL_DFF_X al_c364f203 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[57]));
  AL_DFF_X al_19d3bed2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[58]));
  AL_DFF_X al_f0296ba3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[59]));
  AL_DFF_X al_82a4daff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[60]));
  AL_DFF_X al_88fbc57f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[61]));
  AL_DFF_X al_e66059e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_297c219f[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e95330c[62]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_d0c8e7ec (
    .a(1'b0),
    .o({al_631fb54,open_n32}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3b312457 (
    .a(al_174c5039[32]),
    .b(al_297c219f[32]),
    .c(al_631fb54),
    .o({al_6a2b173c,al_e6544b06[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dd806e4f (
    .a(al_174c5039[33]),
    .b(al_297c219f[33]),
    .c(al_6a2b173c),
    .o({al_c111311e,al_e6544b06[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e3cae714 (
    .a(al_174c5039[34]),
    .b(al_297c219f[34]),
    .c(al_c111311e),
    .o({al_a67d66f1,al_e6544b06[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_21b6413c (
    .a(al_174c5039[35]),
    .b(al_297c219f[35]),
    .c(al_a67d66f1),
    .o({al_5cbcdb58,al_e6544b06[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4828c238 (
    .a(al_174c5039[36]),
    .b(al_297c219f[36]),
    .c(al_5cbcdb58),
    .o({al_bb2c445c,al_e6544b06[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_91cf1d4d (
    .a(al_174c5039[37]),
    .b(al_297c219f[37]),
    .c(al_bb2c445c),
    .o({al_a217d3f1,al_e6544b06[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_65e38deb (
    .a(al_174c5039[38]),
    .b(al_297c219f[38]),
    .c(al_a217d3f1),
    .o({al_5cde9409,al_e6544b06[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c55c685a (
    .a(al_174c5039[39]),
    .b(al_297c219f[39]),
    .c(al_5cde9409),
    .o({al_7b31c923,al_e6544b06[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc86b8ba (
    .a(al_174c5039[40]),
    .b(al_297c219f[40]),
    .c(al_7b31c923),
    .o({al_855bfb89,al_e6544b06[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ac0218f3 (
    .a(al_174c5039[41]),
    .b(al_297c219f[41]),
    .c(al_855bfb89),
    .o({al_c41c8842,al_e6544b06[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_36d78fc (
    .a(al_174c5039[42]),
    .b(al_297c219f[42]),
    .c(al_c41c8842),
    .o({al_29e9ad49,al_e6544b06[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_870f13a3 (
    .a(al_174c5039[43]),
    .b(al_297c219f[43]),
    .c(al_29e9ad49),
    .o({al_786a64be,al_e6544b06[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_61a0d7ee (
    .a(al_174c5039[44]),
    .b(al_297c219f[44]),
    .c(al_786a64be),
    .o({al_9b1b3762,al_e6544b06[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd9c53 (
    .a(al_174c5039[45]),
    .b(al_297c219f[45]),
    .c(al_9b1b3762),
    .o({al_371bfa10,al_e6544b06[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_614e94eb (
    .a(al_174c5039[46]),
    .b(al_297c219f[46]),
    .c(al_371bfa10),
    .o({al_eea0690a,al_e6544b06[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_56056eb (
    .a(al_174c5039[47]),
    .b(al_297c219f[47]),
    .c(al_eea0690a),
    .o({al_670e1d07,al_e6544b06[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_257a444d (
    .c(al_670e1d07),
    .o({open_n35,al_e6544b06[16]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7c262a (
    .a(al_35b24b05),
    .b(al_174c5039[32]),
    .c(al_e6544b06[0]),
    .o(al_45052583[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_272cb0ca (
    .a(al_35b24b05),
    .b(al_174c5039[33]),
    .c(al_e6544b06[1]),
    .o(al_45052583[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4ac007ca (
    .a(al_35b24b05),
    .b(al_174c5039[34]),
    .c(al_e6544b06[2]),
    .o(al_45052583[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b4cbc674 (
    .a(al_35b24b05),
    .b(al_174c5039[35]),
    .c(al_e6544b06[3]),
    .o(al_45052583[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f1b4b396 (
    .a(al_35b24b05),
    .b(al_174c5039[36]),
    .c(al_e6544b06[4]),
    .o(al_45052583[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_67c09b2c (
    .a(al_35b24b05),
    .b(al_174c5039[37]),
    .c(al_e6544b06[5]),
    .o(al_45052583[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5943e37e (
    .a(al_35b24b05),
    .b(al_174c5039[38]),
    .c(al_e6544b06[6]),
    .o(al_45052583[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f4a20a75 (
    .a(al_35b24b05),
    .b(al_174c5039[39]),
    .c(al_e6544b06[7]),
    .o(al_45052583[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_851c2339 (
    .a(al_35b24b05),
    .b(al_174c5039[40]),
    .c(al_e6544b06[8]),
    .o(al_45052583[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c79cfdbf (
    .a(al_35b24b05),
    .b(al_174c5039[41]),
    .c(al_e6544b06[9]),
    .o(al_45052583[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f5969b73 (
    .a(al_35b24b05),
    .b(al_174c5039[42]),
    .c(al_e6544b06[10]),
    .o(al_45052583[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2d1bf9cc (
    .a(al_35b24b05),
    .b(al_174c5039[43]),
    .c(al_e6544b06[11]),
    .o(al_45052583[43]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_6f63c383 (
    .a(al_297c219f[58]),
    .b(al_297c219f[59]),
    .c(al_297c219f[60]),
    .d(al_297c219f[61]),
    .e(al_297c219f[62]),
    .f(al_297c219f[63]),
    .o(al_ee69ef7a));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_a6507f59 (
    .a(al_297c219f[52]),
    .b(al_297c219f[53]),
    .c(al_297c219f[54]),
    .d(al_297c219f[55]),
    .e(al_297c219f[56]),
    .f(al_297c219f[57]),
    .o(al_11e5467d));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_954c18ee (
    .a(al_297c219f[48]),
    .b(al_297c219f[49]),
    .c(al_297c219f[50]),
    .d(al_297c219f[51]),
    .e(al_e6544b06[16]),
    .o(al_3910e4e4));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_9a90cfa2 (
    .a(al_ee69ef7a),
    .b(al_11e5467d),
    .c(al_3910e4e4),
    .o(al_35b24b05));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b925fc76 (
    .a(al_35b24b05),
    .b(al_174c5039[44]),
    .c(al_e6544b06[12]),
    .o(al_45052583[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ee1e7af6 (
    .a(al_35b24b05),
    .b(al_174c5039[45]),
    .c(al_e6544b06[13]),
    .o(al_45052583[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bb58c7b6 (
    .a(al_35b24b05),
    .b(al_174c5039[46]),
    .c(al_e6544b06[14]),
    .o(al_45052583[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f5635f95 (
    .a(al_35b24b05),
    .b(al_174c5039[47]),
    .c(al_e6544b06[15]),
    .o(al_45052583[47]));
  AL_DFF_X al_73d1c90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[0]));
  AL_DFF_X al_387f0ce1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[9]));
  AL_DFF_X al_baeaa68c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[10]));
  AL_DFF_X al_cdb41423 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[11]));
  AL_DFF_X al_8875db47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[12]));
  AL_DFF_X al_3e11e321 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[13]));
  AL_DFF_X al_2c2ab09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[14]));
  AL_DFF_X al_5591d838 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[15]));
  AL_DFF_X al_12a9d470 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[16]));
  AL_DFF_X al_b4675e5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[17]));
  AL_DFF_X al_6d398222 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[18]));
  AL_DFF_X al_c254c362 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[1]));
  AL_DFF_X al_9c3707df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[19]));
  AL_DFF_X al_c1e88f58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[20]));
  AL_DFF_X al_6bbd0477 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[21]));
  AL_DFF_X al_d8a27b85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[22]));
  AL_DFF_X al_b7425df8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[23]));
  AL_DFF_X al_edd1b008 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[24]));
  AL_DFF_X al_7450cf1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[25]));
  AL_DFF_X al_212255eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[26]));
  AL_DFF_X al_71b36ee5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[27]));
  AL_DFF_X al_4a39527f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[28]));
  AL_DFF_X al_78b74f15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[2]));
  AL_DFF_X al_e42f7f42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[29]));
  AL_DFF_X al_ca5de5cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[30]));
  AL_DFF_X al_369be645 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[31]));
  AL_DFF_X al_a1c4afd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[32]));
  AL_DFF_X al_dcf4cd32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[33]));
  AL_DFF_X al_db42196e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[34]));
  AL_DFF_X al_34f25408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[35]));
  AL_DFF_X al_54add82c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[36]));
  AL_DFF_X al_c1a742a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[37]));
  AL_DFF_X al_26b47b2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[38]));
  AL_DFF_X al_173e7559 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[3]));
  AL_DFF_X al_cd9686c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[39]));
  AL_DFF_X al_f3066eec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[40]));
  AL_DFF_X al_fec4ecd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[41]));
  AL_DFF_X al_eb22b23a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[42]));
  AL_DFF_X al_a2cd5af9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[43]));
  AL_DFF_X al_ce580533 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[44]));
  AL_DFF_X al_63c5bbef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[45]));
  AL_DFF_X al_62177e2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[46]));
  AL_DFF_X al_2e6d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_45052583[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[47]));
  AL_DFF_X al_68536e25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[4]));
  AL_DFF_X al_4ecd45f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[5]));
  AL_DFF_X al_cd5f5f4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[6]));
  AL_DFF_X al_e8c12bf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[7]));
  AL_DFF_X al_5adb0590 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_174c5039[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1276f4f7[8]));
  AL_DFF_X al_7fbf5c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35b24b05),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[0]));
  AL_DFF_X al_6f0aaea3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[9]));
  AL_DFF_X al_1ce6b5a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[10]));
  AL_DFF_X al_d9342534 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[11]));
  AL_DFF_X al_c69f5023 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[12]));
  AL_DFF_X al_1e189ba4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[13]));
  AL_DFF_X al_7bde4041 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[14]));
  AL_DFF_X al_7dd6e87e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[15]));
  AL_DFF_X al_aff378f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[1]));
  AL_DFF_X al_d90e47d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[2]));
  AL_DFF_X al_a86140b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[3]));
  AL_DFF_X al_c2e35613 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[4]));
  AL_DFF_X al_c182e813 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[5]));
  AL_DFF_X al_74a46fd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[6]));
  AL_DFF_X al_25697b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[7]));
  AL_DFF_X al_9ac728f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebfa785c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4daf6f3[8]));
  AL_DFF_X al_90b6272a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5ed5f44b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_54284e1f[0]));
  AL_DFF_X al_410157de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[30]));
  AL_DFF_X al_e79c25a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[31]));
  AL_DFF_X al_73b78957 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[32]));
  AL_DFF_X al_a6829b65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[33]));
  AL_DFF_X al_4baad3a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[34]));
  AL_DFF_X al_d262cf0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[35]));
  AL_DFF_X al_f8581787 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[36]));
  AL_DFF_X al_1776b692 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[37]));
  AL_DFF_X al_674e70fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[38]));
  AL_DFF_X al_75d7aff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[39]));
  AL_DFF_X al_22620f95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[40]));
  AL_DFF_X al_26e967a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[41]));
  AL_DFF_X al_71882c8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[42]));
  AL_DFF_X al_b1e7dc15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[43]));
  AL_DFF_X al_600a58e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[44]));
  AL_DFF_X al_49a8d07f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[45]));
  AL_DFF_X al_ef8917f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[46]));
  AL_DFF_X al_38ad3501 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[47]));
  AL_DFF_X al_f9d48560 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[48]));
  AL_DFF_X al_a0df6e34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[49]));
  AL_DFF_X al_c00f4f17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[50]));
  AL_DFF_X al_c9be8077 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[51]));
  AL_DFF_X al_21ed5e97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[52]));
  AL_DFF_X al_986f2199 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[53]));
  AL_DFF_X al_6a2ac330 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[54]));
  AL_DFF_X al_b4987f20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[55]));
  AL_DFF_X al_7c4bcbd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[56]));
  AL_DFF_X al_b6c04ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[57]));
  AL_DFF_X al_e3caa495 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[58]));
  AL_DFF_X al_6208af5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[59]));
  AL_DFF_X al_1d278f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[60]));
  AL_DFF_X al_35996807 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e95330c[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b4e2b23b[61]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_6fcf33ef (
    .a(1'b0),
    .o({al_61d00fc7,open_n38}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1f18f11 (
    .a(al_1276f4f7[31]),
    .b(al_2e95330c[31]),
    .c(al_61d00fc7),
    .o({al_550f60c3,al_eab6bdfe[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2a91fb6a (
    .a(al_1276f4f7[32]),
    .b(al_2e95330c[32]),
    .c(al_550f60c3),
    .o({al_5f55c3b4,al_eab6bdfe[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_262bc5a2 (
    .a(al_1276f4f7[33]),
    .b(al_2e95330c[33]),
    .c(al_5f55c3b4),
    .o({al_dc7a89a9,al_eab6bdfe[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3e6b047a (
    .a(al_1276f4f7[34]),
    .b(al_2e95330c[34]),
    .c(al_dc7a89a9),
    .o({al_5aec0d3d,al_eab6bdfe[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_29fab510 (
    .a(al_1276f4f7[35]),
    .b(al_2e95330c[35]),
    .c(al_5aec0d3d),
    .o({al_146c9954,al_eab6bdfe[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_db23ffd5 (
    .a(al_1276f4f7[36]),
    .b(al_2e95330c[36]),
    .c(al_146c9954),
    .o({al_95294fb6,al_eab6bdfe[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5484049c (
    .a(al_1276f4f7[37]),
    .b(al_2e95330c[37]),
    .c(al_95294fb6),
    .o({al_2b309dfb,al_eab6bdfe[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_428c239c (
    .a(al_1276f4f7[38]),
    .b(al_2e95330c[38]),
    .c(al_2b309dfb),
    .o({al_af8062a0,al_eab6bdfe[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fcbddfe9 (
    .a(al_1276f4f7[39]),
    .b(al_2e95330c[39]),
    .c(al_af8062a0),
    .o({al_3c2e3c3a,al_eab6bdfe[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2611368e (
    .a(al_1276f4f7[40]),
    .b(al_2e95330c[40]),
    .c(al_3c2e3c3a),
    .o({al_b4c76c23,al_eab6bdfe[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f40d993a (
    .a(al_1276f4f7[41]),
    .b(al_2e95330c[41]),
    .c(al_b4c76c23),
    .o({al_bcaace37,al_eab6bdfe[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f2c37936 (
    .a(al_1276f4f7[42]),
    .b(al_2e95330c[42]),
    .c(al_bcaace37),
    .o({al_6dbf3665,al_eab6bdfe[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f8b84eb9 (
    .a(al_1276f4f7[43]),
    .b(al_2e95330c[43]),
    .c(al_6dbf3665),
    .o({al_8a54e775,al_eab6bdfe[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2de59830 (
    .a(al_1276f4f7[44]),
    .b(al_2e95330c[44]),
    .c(al_8a54e775),
    .o({al_8f1f7251,al_eab6bdfe[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d968dd9d (
    .a(al_1276f4f7[45]),
    .b(al_2e95330c[45]),
    .c(al_8f1f7251),
    .o({al_eb782a2a,al_eab6bdfe[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c0bdc2cd (
    .a(al_1276f4f7[46]),
    .b(al_2e95330c[46]),
    .c(al_eb782a2a),
    .o({al_d3a3aa84,al_eab6bdfe[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b3f3da0 (
    .a(al_1276f4f7[47]),
    .b(al_2e95330c[47]),
    .c(al_d3a3aa84),
    .o({al_43acb4d3,al_eab6bdfe[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6eec3940 (
    .c(al_43acb4d3),
    .o({open_n41,al_eab6bdfe[17]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_14a69f62 (
    .a(al_2e95330c[58]),
    .b(al_2e95330c[59]),
    .c(al_2e95330c[60]),
    .d(al_2e95330c[61]),
    .e(al_2e95330c[62]),
    .f(al_eab6bdfe[17]),
    .o(al_2a00900c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_7c78ef94 (
    .a(al_2e95330c[52]),
    .b(al_2e95330c[53]),
    .c(al_2e95330c[54]),
    .d(al_2e95330c[55]),
    .e(al_2e95330c[56]),
    .f(al_2e95330c[57]),
    .o(al_66810f7a));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_d77dde98 (
    .a(al_2a00900c),
    .b(al_66810f7a),
    .c(al_2e95330c[48]),
    .d(al_2e95330c[49]),
    .e(al_2e95330c[50]),
    .f(al_2e95330c[51]),
    .o(al_dbcf415b));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dfedf33e (
    .a(al_dbcf415b),
    .b(al_1276f4f7[31]),
    .c(al_eab6bdfe[0]),
    .o(al_b5df9b8a[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_745c26b7 (
    .a(al_dbcf415b),
    .b(al_1276f4f7[32]),
    .c(al_eab6bdfe[1]),
    .o(al_b5df9b8a[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_927b78fa (
    .a(al_dbcf415b),
    .b(al_1276f4f7[33]),
    .c(al_eab6bdfe[2]),
    .o(al_b5df9b8a[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2bc7c239 (
    .a(al_dbcf415b),
    .b(al_1276f4f7[34]),
    .c(al_eab6bdfe[3]),
    .o(al_b5df9b8a[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fe7d7f2c (
    .a(al_dbcf415b),
    .b(al_1276f4f7[35]),
    .c(al_eab6bdfe[4]),
    .o(al_b5df9b8a[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b4b2ac09 (
    .a(al_dbcf415b),
    .b(al_1276f4f7[36]),
    .c(al_eab6bdfe[5]),
    .o(al_b5df9b8a[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_615d6af (
    .a(al_dbcf415b),
    .b(al_1276f4f7[37]),
    .c(al_eab6bdfe[6]),
    .o(al_b5df9b8a[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_36ce12b0 (
    .a(al_dbcf415b),
    .b(al_1276f4f7[38]),
    .c(al_eab6bdfe[7]),
    .o(al_b5df9b8a[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_48df1a2c (
    .a(al_dbcf415b),
    .b(al_1276f4f7[39]),
    .c(al_eab6bdfe[8]),
    .o(al_b5df9b8a[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_11394d2d (
    .a(al_dbcf415b),
    .b(al_1276f4f7[40]),
    .c(al_eab6bdfe[9]),
    .o(al_b5df9b8a[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bbc02865 (
    .a(al_dbcf415b),
    .b(al_1276f4f7[41]),
    .c(al_eab6bdfe[10]),
    .o(al_b5df9b8a[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1086896d (
    .a(al_dbcf415b),
    .b(al_1276f4f7[42]),
    .c(al_eab6bdfe[11]),
    .o(al_b5df9b8a[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9593cd72 (
    .a(al_dbcf415b),
    .b(al_1276f4f7[43]),
    .c(al_eab6bdfe[12]),
    .o(al_b5df9b8a[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b42d475e (
    .a(al_dbcf415b),
    .b(al_1276f4f7[44]),
    .c(al_eab6bdfe[13]),
    .o(al_b5df9b8a[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_81881895 (
    .a(al_dbcf415b),
    .b(al_1276f4f7[45]),
    .c(al_eab6bdfe[14]),
    .o(al_b5df9b8a[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e702841e (
    .a(al_dbcf415b),
    .b(al_1276f4f7[46]),
    .c(al_eab6bdfe[15]),
    .o(al_b5df9b8a[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6c01d9a3 (
    .a(al_dbcf415b),
    .b(al_1276f4f7[47]),
    .c(al_eab6bdfe[16]),
    .o(al_b5df9b8a[47]));
  AL_DFF_X al_8228c33b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[0]));
  AL_DFF_X al_63689616 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[9]));
  AL_DFF_X al_7b1735a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[10]));
  AL_DFF_X al_7c02935a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[11]));
  AL_DFF_X al_dcda2fe8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[12]));
  AL_DFF_X al_cf1c52ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[13]));
  AL_DFF_X al_8cfeef6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[14]));
  AL_DFF_X al_1123f9aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[15]));
  AL_DFF_X al_25c62528 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[16]));
  AL_DFF_X al_9df6fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[17]));
  AL_DFF_X al_4b822ec3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[18]));
  AL_DFF_X al_38207d0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[1]));
  AL_DFF_X al_21f382b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[19]));
  AL_DFF_X al_8fa02dee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[20]));
  AL_DFF_X al_e0ffb31e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[21]));
  AL_DFF_X al_32673cbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[22]));
  AL_DFF_X al_7970e9a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[23]));
  AL_DFF_X al_140cb0a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[24]));
  AL_DFF_X al_1a038fd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[25]));
  AL_DFF_X al_34873373 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[26]));
  AL_DFF_X al_6124fd4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[27]));
  AL_DFF_X al_8c96d098 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[28]));
  AL_DFF_X al_f8653e31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[2]));
  AL_DFF_X al_d01db61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[29]));
  AL_DFF_X al_d60f399e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[30]));
  AL_DFF_X al_1ff19ca9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[31]));
  AL_DFF_X al_a5eb91f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[32]));
  AL_DFF_X al_a0acc29b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[33]));
  AL_DFF_X al_d6502a1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[34]));
  AL_DFF_X al_36327b43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[35]));
  AL_DFF_X al_3a8a806e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[36]));
  AL_DFF_X al_d8582c9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[37]));
  AL_DFF_X al_c792578d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[38]));
  AL_DFF_X al_f92d7dae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[3]));
  AL_DFF_X al_f7abc49c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[39]));
  AL_DFF_X al_4c6ea502 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[40]));
  AL_DFF_X al_1f928eca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[41]));
  AL_DFF_X al_f6606f85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[42]));
  AL_DFF_X al_8f3e7581 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[43]));
  AL_DFF_X al_9c326d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[44]));
  AL_DFF_X al_128bfd95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[45]));
  AL_DFF_X al_b29e0cf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[46]));
  AL_DFF_X al_b724ce39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b5df9b8a[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[47]));
  AL_DFF_X al_dc910a91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[4]));
  AL_DFF_X al_3e444bb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[5]));
  AL_DFF_X al_561b3b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[6]));
  AL_DFF_X al_a50b8fb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[7]));
  AL_DFF_X al_a0dfbce8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1276f4f7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3692f86e[8]));
  AL_DFF_X al_57f4ea38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dbcf415b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[0]));
  AL_DFF_X al_5df86358 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[9]));
  AL_DFF_X al_64776e57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[10]));
  AL_DFF_X al_10b1ee75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[11]));
  AL_DFF_X al_8ac52804 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[12]));
  AL_DFF_X al_3a300584 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[13]));
  AL_DFF_X al_d39e4391 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[14]));
  AL_DFF_X al_c0df65c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[15]));
  AL_DFF_X al_334e5fcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[16]));
  AL_DFF_X al_a74836b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[1]));
  AL_DFF_X al_e8e7348d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[2]));
  AL_DFF_X al_2d83f6b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[3]));
  AL_DFF_X al_b517c6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[4]));
  AL_DFF_X al_33454ea9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[5]));
  AL_DFF_X al_181dcb10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[6]));
  AL_DFF_X al_8fdb623 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[7]));
  AL_DFF_X al_a8fa6efb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4daf6f3[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c94ca47[8]));
  AL_DFF_X al_3d0e33d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_54284e1f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f83a6cd4[0]));
  AL_DFF_X al_5a175824 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[29]));
  AL_DFF_X al_6ca055de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[30]));
  AL_DFF_X al_8e54175e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[31]));
  AL_DFF_X al_168df569 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[32]));
  AL_DFF_X al_cf731055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[33]));
  AL_DFF_X al_60db824f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[34]));
  AL_DFF_X al_2871124b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[35]));
  AL_DFF_X al_996be600 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[36]));
  AL_DFF_X al_1ecadc14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[37]));
  AL_DFF_X al_74e86b34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[38]));
  AL_DFF_X al_54a99f79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[39]));
  AL_DFF_X al_392b3949 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[40]));
  AL_DFF_X al_da323314 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[41]));
  AL_DFF_X al_9b46d608 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[42]));
  AL_DFF_X al_1fead1c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[43]));
  AL_DFF_X al_d62a8a7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[44]));
  AL_DFF_X al_f40789a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[45]));
  AL_DFF_X al_62bd195f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[46]));
  AL_DFF_X al_50c85c5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[47]));
  AL_DFF_X al_7b612d55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[48]));
  AL_DFF_X al_9a6652cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[49]));
  AL_DFF_X al_5bbf6088 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[50]));
  AL_DFF_X al_111dfb40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[51]));
  AL_DFF_X al_92e20209 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[52]));
  AL_DFF_X al_a594aa6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[53]));
  AL_DFF_X al_8aae83ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[54]));
  AL_DFF_X al_5347786f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[55]));
  AL_DFF_X al_e53b3157 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[56]));
  AL_DFF_X al_78da4828 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[57]));
  AL_DFF_X al_ef297d08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[58]));
  AL_DFF_X al_f4bb89d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[59]));
  AL_DFF_X al_5bd48ed4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b4e2b23b[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7d838f[60]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_18ac468c (
    .a(1'b0),
    .o({al_e40ec610,open_n44}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4accccca (
    .a(al_3692f86e[30]),
    .b(al_b4e2b23b[30]),
    .c(al_e40ec610),
    .o({al_3ca88873,al_7bf458d0[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_250ef0cd (
    .a(al_3692f86e[31]),
    .b(al_b4e2b23b[31]),
    .c(al_3ca88873),
    .o({al_4ff8e4,al_7bf458d0[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_952d8070 (
    .a(al_3692f86e[32]),
    .b(al_b4e2b23b[32]),
    .c(al_4ff8e4),
    .o({al_cd79137f,al_7bf458d0[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7ede1b70 (
    .a(al_3692f86e[33]),
    .b(al_b4e2b23b[33]),
    .c(al_cd79137f),
    .o({al_dbca7fa0,al_7bf458d0[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_20307fd (
    .a(al_3692f86e[34]),
    .b(al_b4e2b23b[34]),
    .c(al_dbca7fa0),
    .o({al_547f2817,al_7bf458d0[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1969127d (
    .a(al_3692f86e[35]),
    .b(al_b4e2b23b[35]),
    .c(al_547f2817),
    .o({al_85dc8a57,al_7bf458d0[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bb7d2346 (
    .a(al_3692f86e[36]),
    .b(al_b4e2b23b[36]),
    .c(al_85dc8a57),
    .o({al_2ed9b6e7,al_7bf458d0[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fe4fc43b (
    .a(al_3692f86e[37]),
    .b(al_b4e2b23b[37]),
    .c(al_2ed9b6e7),
    .o({al_283f9817,al_7bf458d0[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dafd66b5 (
    .a(al_3692f86e[38]),
    .b(al_b4e2b23b[38]),
    .c(al_283f9817),
    .o({al_1967a37e,al_7bf458d0[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4b6f18f2 (
    .a(al_3692f86e[39]),
    .b(al_b4e2b23b[39]),
    .c(al_1967a37e),
    .o({al_32707238,al_7bf458d0[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8e1c57b (
    .a(al_3692f86e[40]),
    .b(al_b4e2b23b[40]),
    .c(al_32707238),
    .o({al_2c79b8f0,al_7bf458d0[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f78e0b95 (
    .a(al_3692f86e[41]),
    .b(al_b4e2b23b[41]),
    .c(al_2c79b8f0),
    .o({al_6fa79631,al_7bf458d0[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_49411112 (
    .a(al_3692f86e[42]),
    .b(al_b4e2b23b[42]),
    .c(al_6fa79631),
    .o({al_683a8463,al_7bf458d0[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4cb6a96c (
    .a(al_3692f86e[43]),
    .b(al_b4e2b23b[43]),
    .c(al_683a8463),
    .o({al_c6efb15f,al_7bf458d0[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6d616ad8 (
    .a(al_3692f86e[44]),
    .b(al_b4e2b23b[44]),
    .c(al_c6efb15f),
    .o({al_16cee9f7,al_7bf458d0[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4d0fc331 (
    .a(al_3692f86e[45]),
    .b(al_b4e2b23b[45]),
    .c(al_16cee9f7),
    .o({al_33147ecd,al_7bf458d0[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6326be7f (
    .a(al_3692f86e[46]),
    .b(al_b4e2b23b[46]),
    .c(al_33147ecd),
    .o({al_7644ebe6,al_7bf458d0[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7f41e945 (
    .a(al_3692f86e[47]),
    .b(al_b4e2b23b[47]),
    .c(al_7644ebe6),
    .o({al_a21a5b9f,al_7bf458d0[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a215114 (
    .c(al_a21a5b9f),
    .o({open_n47,al_7bf458d0[18]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_85f25e31 (
    .a(al_a7eb7389),
    .b(al_3692f86e[30]),
    .c(al_7bf458d0[0]),
    .o(al_28955387[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5542f9f5 (
    .a(al_a7eb7389),
    .b(al_3692f86e[31]),
    .c(al_7bf458d0[1]),
    .o(al_28955387[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_28d9af9e (
    .a(al_a7eb7389),
    .b(al_3692f86e[32]),
    .c(al_7bf458d0[2]),
    .o(al_28955387[32]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_ebf88f57 (
    .a(al_b4e2b23b[56]),
    .b(al_b4e2b23b[57]),
    .c(al_b4e2b23b[58]),
    .d(al_b4e2b23b[59]),
    .e(al_b4e2b23b[60]),
    .f(al_b4e2b23b[61]),
    .o(al_84143d7e));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_b1895f93 (
    .a(al_b4e2b23b[50]),
    .b(al_b4e2b23b[51]),
    .c(al_b4e2b23b[52]),
    .d(al_b4e2b23b[53]),
    .e(al_b4e2b23b[54]),
    .f(al_b4e2b23b[55]),
    .o(al_2e9e4aac));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    al_35278270 (
    .a(al_84143d7e),
    .b(al_2e9e4aac),
    .c(al_b4e2b23b[48]),
    .d(al_b4e2b23b[49]),
    .e(al_7bf458d0[18]),
    .o(al_a7eb7389));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1c1d7f39 (
    .a(al_a7eb7389),
    .b(al_3692f86e[33]),
    .c(al_7bf458d0[3]),
    .o(al_28955387[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a3015a8c (
    .a(al_a7eb7389),
    .b(al_3692f86e[34]),
    .c(al_7bf458d0[4]),
    .o(al_28955387[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ab0a9c45 (
    .a(al_a7eb7389),
    .b(al_3692f86e[35]),
    .c(al_7bf458d0[5]),
    .o(al_28955387[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1e0b59ca (
    .a(al_a7eb7389),
    .b(al_3692f86e[36]),
    .c(al_7bf458d0[6]),
    .o(al_28955387[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_de1c54c (
    .a(al_a7eb7389),
    .b(al_3692f86e[37]),
    .c(al_7bf458d0[7]),
    .o(al_28955387[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_41673ad6 (
    .a(al_a7eb7389),
    .b(al_3692f86e[38]),
    .c(al_7bf458d0[8]),
    .o(al_28955387[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_61bd199a (
    .a(al_a7eb7389),
    .b(al_3692f86e[39]),
    .c(al_7bf458d0[9]),
    .o(al_28955387[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9a0cf1e (
    .a(al_a7eb7389),
    .b(al_3692f86e[40]),
    .c(al_7bf458d0[10]),
    .o(al_28955387[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fcf2e794 (
    .a(al_a7eb7389),
    .b(al_3692f86e[41]),
    .c(al_7bf458d0[11]),
    .o(al_28955387[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_aebdb2bc (
    .a(al_a7eb7389),
    .b(al_3692f86e[42]),
    .c(al_7bf458d0[12]),
    .o(al_28955387[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c9a31461 (
    .a(al_a7eb7389),
    .b(al_3692f86e[43]),
    .c(al_7bf458d0[13]),
    .o(al_28955387[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3a849325 (
    .a(al_a7eb7389),
    .b(al_3692f86e[44]),
    .c(al_7bf458d0[14]),
    .o(al_28955387[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1050c744 (
    .a(al_a7eb7389),
    .b(al_3692f86e[45]),
    .c(al_7bf458d0[15]),
    .o(al_28955387[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_68d574d1 (
    .a(al_a7eb7389),
    .b(al_3692f86e[46]),
    .c(al_7bf458d0[16]),
    .o(al_28955387[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a1c84e69 (
    .a(al_a7eb7389),
    .b(al_3692f86e[47]),
    .c(al_7bf458d0[17]),
    .o(al_28955387[47]));
  AL_DFF_X al_18bb1de8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[0]));
  AL_DFF_X al_776d3244 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[9]));
  AL_DFF_X al_d53f9762 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[10]));
  AL_DFF_X al_e17dc1af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[11]));
  AL_DFF_X al_a7eb85de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[12]));
  AL_DFF_X al_ad2fe98f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[13]));
  AL_DFF_X al_bf50e8f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[14]));
  AL_DFF_X al_b1791ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[15]));
  AL_DFF_X al_ab996acc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[16]));
  AL_DFF_X al_5c40808e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[17]));
  AL_DFF_X al_4bd7ef6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[18]));
  AL_DFF_X al_a9ab99e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[1]));
  AL_DFF_X al_afb234a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[19]));
  AL_DFF_X al_bd319407 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[20]));
  AL_DFF_X al_674890e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[21]));
  AL_DFF_X al_e4fbd537 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[22]));
  AL_DFF_X al_91552b0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[23]));
  AL_DFF_X al_c3fbc2d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[24]));
  AL_DFF_X al_ca6bab7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[25]));
  AL_DFF_X al_31a6d3c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[26]));
  AL_DFF_X al_4d3464af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[27]));
  AL_DFF_X al_18b33cba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[28]));
  AL_DFF_X al_c3eb797b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[2]));
  AL_DFF_X al_2398c0f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[29]));
  AL_DFF_X al_10f2eddb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[30]));
  AL_DFF_X al_b114c8eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[31]));
  AL_DFF_X al_5b701e40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[32]));
  AL_DFF_X al_d369e009 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[33]));
  AL_DFF_X al_2628ce0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[34]));
  AL_DFF_X al_b04b8988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[35]));
  AL_DFF_X al_dcf44a77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[36]));
  AL_DFF_X al_13ef90c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[37]));
  AL_DFF_X al_6aca39cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[38]));
  AL_DFF_X al_c818e8eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[3]));
  AL_DFF_X al_92350570 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[39]));
  AL_DFF_X al_5f8779f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[40]));
  AL_DFF_X al_dbcf4284 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[41]));
  AL_DFF_X al_231fd662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[42]));
  AL_DFF_X al_b85de882 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[43]));
  AL_DFF_X al_4a5b6b50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[44]));
  AL_DFF_X al_b9e26e55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[45]));
  AL_DFF_X al_a017c387 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[46]));
  AL_DFF_X al_f0ff499f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28955387[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[47]));
  AL_DFF_X al_8d086ce4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[4]));
  AL_DFF_X al_d812c3d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[5]));
  AL_DFF_X al_3aa3fcfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[6]));
  AL_DFF_X al_37c546ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[7]));
  AL_DFF_X al_5e6a990f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3692f86e[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_368cfa5b[8]));
  AL_DFF_X al_1d20e79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a7eb7389),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[0]));
  AL_DFF_X al_db7fb1be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[9]));
  AL_DFF_X al_81a25b86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[10]));
  AL_DFF_X al_f94d695c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[11]));
  AL_DFF_X al_cc2aab77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[12]));
  AL_DFF_X al_fddb39a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[13]));
  AL_DFF_X al_81438fd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[14]));
  AL_DFF_X al_ce956221 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[15]));
  AL_DFF_X al_7a5b7d3d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[16]));
  AL_DFF_X al_ed172cd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[17]));
  AL_DFF_X al_368dd9e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[1]));
  AL_DFF_X al_992a2abb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[2]));
  AL_DFF_X al_348dfd59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[3]));
  AL_DFF_X al_bd3dea9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[4]));
  AL_DFF_X al_44bbf870 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[5]));
  AL_DFF_X al_d9ead8a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[6]));
  AL_DFF_X al_855a5ce3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[7]));
  AL_DFF_X al_4fdb8b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c94ca47[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_def6d145[8]));
  AL_DFF_X al_ed0a0726 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f83a6cd4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b0a2efb7[0]));
  AL_DFF_X al_42678e11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[28]));
  AL_DFF_X al_8530090f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[29]));
  AL_DFF_X al_847212c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[30]));
  AL_DFF_X al_f6faa66c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[31]));
  AL_DFF_X al_21e73ae6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[32]));
  AL_DFF_X al_316c0068 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[33]));
  AL_DFF_X al_9e567d9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[34]));
  AL_DFF_X al_6ab6e965 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[35]));
  AL_DFF_X al_81ee7e6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[36]));
  AL_DFF_X al_413b9952 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[37]));
  AL_DFF_X al_2e676f50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[38]));
  AL_DFF_X al_ade543a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[39]));
  AL_DFF_X al_8db07b94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[40]));
  AL_DFF_X al_3a155b72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[41]));
  AL_DFF_X al_f27218ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[42]));
  AL_DFF_X al_f6fae6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[43]));
  AL_DFF_X al_9f4fee80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[44]));
  AL_DFF_X al_907d37dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[45]));
  AL_DFF_X al_39b523ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[46]));
  AL_DFF_X al_7dbd8a4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[47]));
  AL_DFF_X al_609128e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[48]));
  AL_DFF_X al_fa8bf24f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[49]));
  AL_DFF_X al_14e3a91d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[50]));
  AL_DFF_X al_9aef722f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[51]));
  AL_DFF_X al_28191835 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[52]));
  AL_DFF_X al_1b826c12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[53]));
  AL_DFF_X al_a31f1a8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[54]));
  AL_DFF_X al_1dbd3554 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[55]));
  AL_DFF_X al_ea7465bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[56]));
  AL_DFF_X al_ed329354 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[57]));
  AL_DFF_X al_9a4125e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[58]));
  AL_DFF_X al_7d94eccb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7d838f[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30e951fe[59]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_cda7a94e (
    .a(1'b0),
    .o({al_122ce731,open_n50}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d52d2612 (
    .a(al_368cfa5b[29]),
    .b(al_e7d838f[29]),
    .c(al_122ce731),
    .o({al_93a235f1,al_402e9e3e[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ed2aec00 (
    .a(al_368cfa5b[30]),
    .b(al_e7d838f[30]),
    .c(al_93a235f1),
    .o({al_bfc9143c,al_402e9e3e[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e491932f (
    .a(al_368cfa5b[31]),
    .b(al_e7d838f[31]),
    .c(al_bfc9143c),
    .o({al_8e30be98,al_402e9e3e[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_be22bc88 (
    .a(al_368cfa5b[32]),
    .b(al_e7d838f[32]),
    .c(al_8e30be98),
    .o({al_2ee33b11,al_402e9e3e[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fa37b0ba (
    .a(al_368cfa5b[33]),
    .b(al_e7d838f[33]),
    .c(al_2ee33b11),
    .o({al_cc4f6241,al_402e9e3e[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7546132a (
    .a(al_368cfa5b[34]),
    .b(al_e7d838f[34]),
    .c(al_cc4f6241),
    .o({al_27369a88,al_402e9e3e[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2d94d7aa (
    .a(al_368cfa5b[35]),
    .b(al_e7d838f[35]),
    .c(al_27369a88),
    .o({al_790961ba,al_402e9e3e[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ce58fca0 (
    .a(al_368cfa5b[36]),
    .b(al_e7d838f[36]),
    .c(al_790961ba),
    .o({al_ed8719fc,al_402e9e3e[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c2ef469d (
    .a(al_368cfa5b[37]),
    .b(al_e7d838f[37]),
    .c(al_ed8719fc),
    .o({al_21a14027,al_402e9e3e[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bcd91d6a (
    .a(al_368cfa5b[38]),
    .b(al_e7d838f[38]),
    .c(al_21a14027),
    .o({al_f719f95a,al_402e9e3e[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d058bfd6 (
    .a(al_368cfa5b[39]),
    .b(al_e7d838f[39]),
    .c(al_f719f95a),
    .o({al_eb9006e0,al_402e9e3e[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e5152da0 (
    .a(al_368cfa5b[40]),
    .b(al_e7d838f[40]),
    .c(al_eb9006e0),
    .o({al_6680c576,al_402e9e3e[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9fcb82d8 (
    .a(al_368cfa5b[41]),
    .b(al_e7d838f[41]),
    .c(al_6680c576),
    .o({al_7820cd3f,al_402e9e3e[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_746b42dd (
    .a(al_368cfa5b[42]),
    .b(al_e7d838f[42]),
    .c(al_7820cd3f),
    .o({al_91e67405,al_402e9e3e[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_98ab07dc (
    .a(al_368cfa5b[43]),
    .b(al_e7d838f[43]),
    .c(al_91e67405),
    .o({al_1f539415,al_402e9e3e[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_26555348 (
    .a(al_368cfa5b[44]),
    .b(al_e7d838f[44]),
    .c(al_1f539415),
    .o({al_fdf27789,al_402e9e3e[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4b3a6a81 (
    .a(al_368cfa5b[45]),
    .b(al_e7d838f[45]),
    .c(al_fdf27789),
    .o({al_cd1eb597,al_402e9e3e[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_72a4125e (
    .a(al_368cfa5b[46]),
    .b(al_e7d838f[46]),
    .c(al_cd1eb597),
    .o({al_95c541ba,al_402e9e3e[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a05a31c0 (
    .a(al_368cfa5b[47]),
    .b(al_e7d838f[47]),
    .c(al_95c541ba),
    .o({al_c62ed6f3,al_402e9e3e[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ed6e8571 (
    .c(al_c62ed6f3),
    .o({open_n53,al_402e9e3e[19]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b14aa975 (
    .a(al_3db819db),
    .b(al_368cfa5b[29]),
    .c(al_402e9e3e[0]),
    .o(al_e55e130b[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ee3a7ce4 (
    .a(al_3db819db),
    .b(al_368cfa5b[30]),
    .c(al_402e9e3e[1]),
    .o(al_e55e130b[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f2b14a41 (
    .a(al_3db819db),
    .b(al_368cfa5b[31]),
    .c(al_402e9e3e[2]),
    .o(al_e55e130b[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cbcb2e47 (
    .a(al_3db819db),
    .b(al_368cfa5b[32]),
    .c(al_402e9e3e[3]),
    .o(al_e55e130b[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dba72098 (
    .a(al_3db819db),
    .b(al_368cfa5b[33]),
    .c(al_402e9e3e[4]),
    .o(al_e55e130b[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5a3b106a (
    .a(al_3db819db),
    .b(al_368cfa5b[34]),
    .c(al_402e9e3e[5]),
    .o(al_e55e130b[34]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_eac2ec17 (
    .a(al_e7d838f[56]),
    .b(al_e7d838f[57]),
    .c(al_e7d838f[58]),
    .d(al_e7d838f[59]),
    .e(al_e7d838f[60]),
    .f(al_402e9e3e[19]),
    .o(al_2e458e8c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_2620f3a2 (
    .a(al_e7d838f[50]),
    .b(al_e7d838f[51]),
    .c(al_e7d838f[52]),
    .d(al_e7d838f[53]),
    .e(al_e7d838f[54]),
    .f(al_e7d838f[55]),
    .o(al_314816f3));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_27acf8a6 (
    .a(al_2e458e8c),
    .b(al_314816f3),
    .c(al_e7d838f[48]),
    .d(al_e7d838f[49]),
    .o(al_3db819db));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9af12d8d (
    .a(al_3db819db),
    .b(al_368cfa5b[35]),
    .c(al_402e9e3e[6]),
    .o(al_e55e130b[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8b7adcc5 (
    .a(al_3db819db),
    .b(al_368cfa5b[36]),
    .c(al_402e9e3e[7]),
    .o(al_e55e130b[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a35cdc65 (
    .a(al_3db819db),
    .b(al_368cfa5b[37]),
    .c(al_402e9e3e[8]),
    .o(al_e55e130b[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c4b811e0 (
    .a(al_3db819db),
    .b(al_368cfa5b[38]),
    .c(al_402e9e3e[9]),
    .o(al_e55e130b[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ed727791 (
    .a(al_3db819db),
    .b(al_368cfa5b[39]),
    .c(al_402e9e3e[10]),
    .o(al_e55e130b[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ad81e577 (
    .a(al_3db819db),
    .b(al_368cfa5b[40]),
    .c(al_402e9e3e[11]),
    .o(al_e55e130b[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8631a928 (
    .a(al_3db819db),
    .b(al_368cfa5b[41]),
    .c(al_402e9e3e[12]),
    .o(al_e55e130b[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d48d5725 (
    .a(al_3db819db),
    .b(al_368cfa5b[42]),
    .c(al_402e9e3e[13]),
    .o(al_e55e130b[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_919e35f5 (
    .a(al_3db819db),
    .b(al_368cfa5b[43]),
    .c(al_402e9e3e[14]),
    .o(al_e55e130b[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7ac7f242 (
    .a(al_3db819db),
    .b(al_368cfa5b[44]),
    .c(al_402e9e3e[15]),
    .o(al_e55e130b[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_950b90a1 (
    .a(al_3db819db),
    .b(al_368cfa5b[45]),
    .c(al_402e9e3e[16]),
    .o(al_e55e130b[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_aa784f8c (
    .a(al_3db819db),
    .b(al_368cfa5b[46]),
    .c(al_402e9e3e[17]),
    .o(al_e55e130b[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_718ee93a (
    .a(al_3db819db),
    .b(al_368cfa5b[47]),
    .c(al_402e9e3e[18]),
    .o(al_e55e130b[47]));
  AL_DFF_X al_825b94ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[0]));
  AL_DFF_X al_64686ec5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[9]));
  AL_DFF_X al_c42b06f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[10]));
  AL_DFF_X al_949117cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[11]));
  AL_DFF_X al_b5e1c2a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[12]));
  AL_DFF_X al_b7a26d3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[13]));
  AL_DFF_X al_85170e41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[14]));
  AL_DFF_X al_a733340c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[15]));
  AL_DFF_X al_7590cbf9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[16]));
  AL_DFF_X al_485f20da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[17]));
  AL_DFF_X al_b41efffb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[18]));
  AL_DFF_X al_6a4856ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[1]));
  AL_DFF_X al_6d2b5328 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[19]));
  AL_DFF_X al_7c271034 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[20]));
  AL_DFF_X al_c4131e72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[21]));
  AL_DFF_X al_c7d41878 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[22]));
  AL_DFF_X al_bfad2360 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[23]));
  AL_DFF_X al_f6aace57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[24]));
  AL_DFF_X al_2e9654c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[25]));
  AL_DFF_X al_e3023aa9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[26]));
  AL_DFF_X al_dd645ef2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[27]));
  AL_DFF_X al_b0d35d39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[28]));
  AL_DFF_X al_b9b2e849 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[2]));
  AL_DFF_X al_672e4243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[29]));
  AL_DFF_X al_3b184ac8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[30]));
  AL_DFF_X al_7ab98c24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[31]));
  AL_DFF_X al_d7497b9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[32]));
  AL_DFF_X al_6ed757d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[33]));
  AL_DFF_X al_fd19b0b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[34]));
  AL_DFF_X al_9eeb8748 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[35]));
  AL_DFF_X al_f9321096 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[36]));
  AL_DFF_X al_848e3f39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[37]));
  AL_DFF_X al_a4170a12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[38]));
  AL_DFF_X al_b9f9b6a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[3]));
  AL_DFF_X al_e4a54429 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[39]));
  AL_DFF_X al_437c7fbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[40]));
  AL_DFF_X al_b770a26f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[41]));
  AL_DFF_X al_ba09e6d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[42]));
  AL_DFF_X al_c1a3a539 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[43]));
  AL_DFF_X al_fd6ff08d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[44]));
  AL_DFF_X al_b45a5ce7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[45]));
  AL_DFF_X al_26ec0db0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[46]));
  AL_DFF_X al_1409c98a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e55e130b[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[47]));
  AL_DFF_X al_de3e9208 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[4]));
  AL_DFF_X al_9e981647 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[5]));
  AL_DFF_X al_5a7225d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[6]));
  AL_DFF_X al_39d70248 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[7]));
  AL_DFF_X al_8da03619 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_368cfa5b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e240f99f[8]));
  AL_DFF_X al_1ce013c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3db819db),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[0]));
  AL_DFF_X al_91ba19a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[9]));
  AL_DFF_X al_439e2cf9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[10]));
  AL_DFF_X al_1bbc1fc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[11]));
  AL_DFF_X al_1e26952d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[12]));
  AL_DFF_X al_9b1791be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[13]));
  AL_DFF_X al_e4a1607e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[14]));
  AL_DFF_X al_1953482d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[15]));
  AL_DFF_X al_23b2bef2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[16]));
  AL_DFF_X al_5f4d805e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[17]));
  AL_DFF_X al_6a7e08f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[18]));
  AL_DFF_X al_e785a729 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[1]));
  AL_DFF_X al_949bd746 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[2]));
  AL_DFF_X al_86ad762c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[3]));
  AL_DFF_X al_3398708b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[4]));
  AL_DFF_X al_13d3c4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[5]));
  AL_DFF_X al_94e10038 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[6]));
  AL_DFF_X al_f061bb0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[7]));
  AL_DFF_X al_c311a036 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_def6d145[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf1e6610[8]));
  AL_DFF_X al_2997413d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b0a2efb7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1c8da1e8[0]));
  AL_DFF_X al_705b9202 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[27]));
  AL_DFF_X al_5c0587d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[28]));
  AL_DFF_X al_78960dc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[29]));
  AL_DFF_X al_11ffd508 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[30]));
  AL_DFF_X al_ff127dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[31]));
  AL_DFF_X al_9911ae61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[32]));
  AL_DFF_X al_432689ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[33]));
  AL_DFF_X al_1b945694 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[34]));
  AL_DFF_X al_e98a7f1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[35]));
  AL_DFF_X al_8039622d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[36]));
  AL_DFF_X al_432df7bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[37]));
  AL_DFF_X al_5b978803 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[38]));
  AL_DFF_X al_df7b73b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[39]));
  AL_DFF_X al_5328d756 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[40]));
  AL_DFF_X al_332b1309 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[41]));
  AL_DFF_X al_3e1ee48e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[42]));
  AL_DFF_X al_3d711eb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[43]));
  AL_DFF_X al_8f94578b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[44]));
  AL_DFF_X al_92f4bdaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[45]));
  AL_DFF_X al_ceb3915a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[46]));
  AL_DFF_X al_ad7890f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[47]));
  AL_DFF_X al_e027b850 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[48]));
  AL_DFF_X al_6d101b83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[49]));
  AL_DFF_X al_bca59625 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[50]));
  AL_DFF_X al_19202bca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[51]));
  AL_DFF_X al_1da45e3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[52]));
  AL_DFF_X al_2005ed8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[53]));
  AL_DFF_X al_e37284f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[54]));
  AL_DFF_X al_7056cabd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[55]));
  AL_DFF_X al_22da8370 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[56]));
  AL_DFF_X al_489acad8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[57]));
  AL_DFF_X al_14faedc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30e951fe[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e803eabe[58]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_25b7fcf7 (
    .a(1'b0),
    .o({al_4cb58e58,open_n56}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_52dda05d (
    .a(al_e240f99f[28]),
    .b(al_30e951fe[28]),
    .c(al_4cb58e58),
    .o({al_61f7300c,al_c49873a4[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_24847733 (
    .a(al_e240f99f[29]),
    .b(al_30e951fe[29]),
    .c(al_61f7300c),
    .o({al_51cbf969,al_c49873a4[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c36b179 (
    .a(al_e240f99f[30]),
    .b(al_30e951fe[30]),
    .c(al_51cbf969),
    .o({al_31d377e1,al_c49873a4[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4c002976 (
    .a(al_e240f99f[31]),
    .b(al_30e951fe[31]),
    .c(al_31d377e1),
    .o({al_5e3c7f1a,al_c49873a4[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_350b87d4 (
    .a(al_e240f99f[32]),
    .b(al_30e951fe[32]),
    .c(al_5e3c7f1a),
    .o({al_67c30993,al_c49873a4[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6c41b44d (
    .a(al_e240f99f[33]),
    .b(al_30e951fe[33]),
    .c(al_67c30993),
    .o({al_1c99d5f6,al_c49873a4[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4595b8bb (
    .a(al_e240f99f[34]),
    .b(al_30e951fe[34]),
    .c(al_1c99d5f6),
    .o({al_66df73c7,al_c49873a4[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3867742b (
    .a(al_e240f99f[35]),
    .b(al_30e951fe[35]),
    .c(al_66df73c7),
    .o({al_a3e63ee7,al_c49873a4[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_35e64262 (
    .a(al_e240f99f[36]),
    .b(al_30e951fe[36]),
    .c(al_a3e63ee7),
    .o({al_63d267c1,al_c49873a4[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6fcb7ce (
    .a(al_e240f99f[37]),
    .b(al_30e951fe[37]),
    .c(al_63d267c1),
    .o({al_8aa456b9,al_c49873a4[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b323728 (
    .a(al_e240f99f[38]),
    .b(al_30e951fe[38]),
    .c(al_8aa456b9),
    .o({al_7fa59108,al_c49873a4[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40133431 (
    .a(al_e240f99f[39]),
    .b(al_30e951fe[39]),
    .c(al_7fa59108),
    .o({al_54c1a264,al_c49873a4[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a87c6d02 (
    .a(al_e240f99f[40]),
    .b(al_30e951fe[40]),
    .c(al_54c1a264),
    .o({al_1937c3b1,al_c49873a4[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d1744eaa (
    .a(al_e240f99f[41]),
    .b(al_30e951fe[41]),
    .c(al_1937c3b1),
    .o({al_8d689511,al_c49873a4[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ca1bcb95 (
    .a(al_e240f99f[42]),
    .b(al_30e951fe[42]),
    .c(al_8d689511),
    .o({al_24deb4a,al_c49873a4[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7bf90ede (
    .a(al_e240f99f[43]),
    .b(al_30e951fe[43]),
    .c(al_24deb4a),
    .o({al_38e8d651,al_c49873a4[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9642b13d (
    .a(al_e240f99f[44]),
    .b(al_30e951fe[44]),
    .c(al_38e8d651),
    .o({al_456aad79,al_c49873a4[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8af1f2dd (
    .a(al_e240f99f[45]),
    .b(al_30e951fe[45]),
    .c(al_456aad79),
    .o({al_26b2c4d9,al_c49873a4[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eee40ad9 (
    .a(al_e240f99f[46]),
    .b(al_30e951fe[46]),
    .c(al_26b2c4d9),
    .o({al_9780212c,al_c49873a4[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_de1895e1 (
    .a(al_e240f99f[47]),
    .b(al_30e951fe[47]),
    .c(al_9780212c),
    .o({al_93d510f7,al_c49873a4[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9dc4dee5 (
    .c(al_93d510f7),
    .o({open_n59,al_c49873a4[20]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_862f1392 (
    .a(al_e8916352),
    .b(al_e240f99f[28]),
    .c(al_c49873a4[0]),
    .o(al_abd7cd63[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_165c84e4 (
    .a(al_e8916352),
    .b(al_e240f99f[29]),
    .c(al_c49873a4[1]),
    .o(al_abd7cd63[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dc5f0eed (
    .a(al_e8916352),
    .b(al_e240f99f[30]),
    .c(al_c49873a4[2]),
    .o(al_abd7cd63[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f068bf18 (
    .a(al_e8916352),
    .b(al_e240f99f[31]),
    .c(al_c49873a4[3]),
    .o(al_abd7cd63[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9ce9a74f (
    .a(al_e8916352),
    .b(al_e240f99f[32]),
    .c(al_c49873a4[4]),
    .o(al_abd7cd63[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_97c41c2b (
    .a(al_e8916352),
    .b(al_e240f99f[33]),
    .c(al_c49873a4[5]),
    .o(al_abd7cd63[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d2f70b95 (
    .a(al_e8916352),
    .b(al_e240f99f[34]),
    .c(al_c49873a4[6]),
    .o(al_abd7cd63[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_99ab91f (
    .a(al_e8916352),
    .b(al_e240f99f[35]),
    .c(al_c49873a4[7]),
    .o(al_abd7cd63[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_973f444f (
    .a(al_e8916352),
    .b(al_e240f99f[36]),
    .c(al_c49873a4[8]),
    .o(al_abd7cd63[36]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_55d086f0 (
    .a(al_30e951fe[54]),
    .b(al_30e951fe[55]),
    .c(al_30e951fe[56]),
    .d(al_30e951fe[57]),
    .e(al_30e951fe[58]),
    .f(al_30e951fe[59]),
    .o(al_7cbeb255));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_e72881ef (
    .a(al_30e951fe[48]),
    .b(al_30e951fe[49]),
    .c(al_30e951fe[50]),
    .d(al_30e951fe[51]),
    .e(al_30e951fe[52]),
    .f(al_30e951fe[53]),
    .o(al_5303c8c4));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    al_a4e2475d (
    .a(al_7cbeb255),
    .b(al_5303c8c4),
    .c(al_c49873a4[20]),
    .o(al_e8916352));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3556ea22 (
    .a(al_e8916352),
    .b(al_e240f99f[37]),
    .c(al_c49873a4[9]),
    .o(al_abd7cd63[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_724f15a0 (
    .a(al_e8916352),
    .b(al_e240f99f[38]),
    .c(al_c49873a4[10]),
    .o(al_abd7cd63[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_530c7813 (
    .a(al_e8916352),
    .b(al_e240f99f[39]),
    .c(al_c49873a4[11]),
    .o(al_abd7cd63[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ec1a062f (
    .a(al_e8916352),
    .b(al_e240f99f[40]),
    .c(al_c49873a4[12]),
    .o(al_abd7cd63[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c925d573 (
    .a(al_e8916352),
    .b(al_e240f99f[41]),
    .c(al_c49873a4[13]),
    .o(al_abd7cd63[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e2334a9 (
    .a(al_e8916352),
    .b(al_e240f99f[42]),
    .c(al_c49873a4[14]),
    .o(al_abd7cd63[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9f830702 (
    .a(al_e8916352),
    .b(al_e240f99f[43]),
    .c(al_c49873a4[15]),
    .o(al_abd7cd63[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e8571312 (
    .a(al_e8916352),
    .b(al_e240f99f[44]),
    .c(al_c49873a4[16]),
    .o(al_abd7cd63[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d278ccec (
    .a(al_e8916352),
    .b(al_e240f99f[45]),
    .c(al_c49873a4[17]),
    .o(al_abd7cd63[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_90237383 (
    .a(al_e8916352),
    .b(al_e240f99f[46]),
    .c(al_c49873a4[18]),
    .o(al_abd7cd63[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_29be8fed (
    .a(al_e8916352),
    .b(al_e240f99f[47]),
    .c(al_c49873a4[19]),
    .o(al_abd7cd63[47]));
  AL_DFF_X al_faeae7d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[0]));
  AL_DFF_X al_62d986a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[9]));
  AL_DFF_X al_f5ab8379 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[10]));
  AL_DFF_X al_63a32662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[11]));
  AL_DFF_X al_caf85032 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[12]));
  AL_DFF_X al_1040159e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[13]));
  AL_DFF_X al_94c81132 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[14]));
  AL_DFF_X al_b2ac6d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[15]));
  AL_DFF_X al_33dc707f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[16]));
  AL_DFF_X al_52a56979 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[17]));
  AL_DFF_X al_e572f052 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[18]));
  AL_DFF_X al_e9a04d34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[1]));
  AL_DFF_X al_f0f18f8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[19]));
  AL_DFF_X al_a5c83d1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[20]));
  AL_DFF_X al_ddcc0253 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[21]));
  AL_DFF_X al_c30eda18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[22]));
  AL_DFF_X al_7858d879 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[23]));
  AL_DFF_X al_c4ae18f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[24]));
  AL_DFF_X al_b85c8ede (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[25]));
  AL_DFF_X al_7d39c1de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[26]));
  AL_DFF_X al_c065d63d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[27]));
  AL_DFF_X al_f059b5f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[28]));
  AL_DFF_X al_f311b755 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[2]));
  AL_DFF_X al_c6659043 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[29]));
  AL_DFF_X al_142b4c81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[30]));
  AL_DFF_X al_30a301a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[31]));
  AL_DFF_X al_89db565b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[32]));
  AL_DFF_X al_7cf5596d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[33]));
  AL_DFF_X al_338afd09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[34]));
  AL_DFF_X al_c07a856 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[35]));
  AL_DFF_X al_a100390a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[36]));
  AL_DFF_X al_7b8e0970 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[37]));
  AL_DFF_X al_3a6bb9f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[38]));
  AL_DFF_X al_a1ae0594 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[3]));
  AL_DFF_X al_ae85971f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[39]));
  AL_DFF_X al_af9ecdb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[40]));
  AL_DFF_X al_1eb1dd2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[41]));
  AL_DFF_X al_ccc251e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[42]));
  AL_DFF_X al_1e73c49c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[43]));
  AL_DFF_X al_d3c3306f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[44]));
  AL_DFF_X al_96755eab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[45]));
  AL_DFF_X al_ab691d77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[46]));
  AL_DFF_X al_8b7ba30d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_abd7cd63[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[47]));
  AL_DFF_X al_7ff32e5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[4]));
  AL_DFF_X al_d8a1706f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[5]));
  AL_DFF_X al_35794404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[6]));
  AL_DFF_X al_6a527a68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[7]));
  AL_DFF_X al_af62df4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e240f99f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_80a0f09e[8]));
  AL_DFF_X al_d5f6ba4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e8916352),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[0]));
  AL_DFF_X al_ea4d0f5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[9]));
  AL_DFF_X al_2d20d0c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[10]));
  AL_DFF_X al_4632f197 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[11]));
  AL_DFF_X al_46ac4a06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[12]));
  AL_DFF_X al_9f75d222 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[13]));
  AL_DFF_X al_f62ed231 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[14]));
  AL_DFF_X al_3b6bdbb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[15]));
  AL_DFF_X al_f4aef84c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[16]));
  AL_DFF_X al_7c95736b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[17]));
  AL_DFF_X al_c4e732e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[18]));
  AL_DFF_X al_7707a88f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[1]));
  AL_DFF_X al_5ca3802e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[19]));
  AL_DFF_X al_9f1f21af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[2]));
  AL_DFF_X al_da6a1dc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[3]));
  AL_DFF_X al_562026da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[4]));
  AL_DFF_X al_8755b9f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[5]));
  AL_DFF_X al_24d02d78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[6]));
  AL_DFF_X al_58343e42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[7]));
  AL_DFF_X al_57e97465 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf1e6610[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bd7f7f17[8]));
  AL_DFF_X al_d95ebc9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3da4ff6f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_67f5b0b3[0]));
  AL_DFF_X al_20442dbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[45]));
  AL_DFF_X al_efd17f14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[46]));
  AL_DFF_X al_3f0986c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[47]));
  AL_DFF_X al_cfb977b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[48]));
  AL_DFF_X al_d2aabb97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[49]));
  AL_DFF_X al_4467f980 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[50]));
  AL_DFF_X al_63e84ddc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[51]));
  AL_DFF_X al_d65237c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[52]));
  AL_DFF_X al_6e2eaf21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[53]));
  AL_DFF_X al_6d2caac5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[54]));
  AL_DFF_X al_8c614a0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[55]));
  AL_DFF_X al_df76a933 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[56]));
  AL_DFF_X al_90c94c47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[57]));
  AL_DFF_X al_6b5b892f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[58]));
  AL_DFF_X al_4f8cfc91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[59]));
  AL_DFF_X al_df679ddb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[60]));
  AL_DFF_X al_552c7f75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[61]));
  AL_DFF_X al_dee96dab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[62]));
  AL_DFF_X al_11d581f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[63]));
  AL_DFF_X al_b2d8b26d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[64]));
  AL_DFF_X al_36fd5654 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[65]));
  AL_DFF_X al_bdb38a43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[66]));
  AL_DFF_X al_a46c3591 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[67]));
  AL_DFF_X al_46d09611 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[68]));
  AL_DFF_X al_3d623382 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[69]));
  AL_DFF_X al_947b31e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[70]));
  AL_DFF_X al_7c52a28a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[71]));
  AL_DFF_X al_ab7ea5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[72]));
  AL_DFF_X al_e0b8ad8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[73]));
  AL_DFF_X al_c98ef919 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[74]));
  AL_DFF_X al_24af8f47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[75]));
  AL_DFF_X al_4b704f0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3bd314e4[77]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a637a32[76]));
  AL_MAP_LUT6 #(
    .EQN("(B*A*(~(D)*~((~E*C))*~(F)+~(D)*~((~E*C))*F+D*~((~E*C))*F+~(D)*(~E*C)*F))"),
    .INIT(64'h8888088800880008))
    al_22a7690c (
    .a(al_3b0f07fc),
    .b(al_fd5ea84d),
    .c(al_3bd314e4[46]),
    .d(al_3bd314e4[47]),
    .e(al_83a08f3f[46]),
    .f(al_83a08f3f[47]),
    .o(al_ff28a985));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_a109ae5b (
    .a(al_3bd314e4[66]),
    .b(al_3bd314e4[69]),
    .c(al_3bd314e4[70]),
    .d(al_3bd314e4[73]),
    .e(al_3bd314e4[75]),
    .f(al_3bd314e4[76]),
    .o(al_1634b160));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    al_3490d663 (
    .a(al_45fda30c),
    .b(al_ca8a5a31),
    .c(al_3bd314e4[51]),
    .d(al_3bd314e4[52]),
    .o(al_fd5ea84d));
  AL_MAP_LUT6 #(
    .EQN("(~((C*B*A))*~(D)*E*~(F)+~((C*B*A))*D*E*~(F)+(C*B*A)*D*E*~(F)+(C*B*A)*~(D)*~(E)*F+~((C*B*A))*~(D)*E*F+~((C*B*A))*D*E*F)"),
    .INIT(64'h7f7f0080ff7f0000))
    al_d1ee308f (
    .a(al_3b0f07fc),
    .b(al_fd5ea84d),
    .c(al_3bd314e4[46]),
    .d(al_3bd314e4[47]),
    .e(al_83a08f3f[46]),
    .f(al_83a08f3f[47]),
    .o(al_89f2771a[46]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_6363a9db (
    .a(al_3bd314e4[55]),
    .b(al_3bd314e4[56]),
    .c(al_3bd314e4[58]),
    .d(al_3bd314e4[61]),
    .e(al_3bd314e4[63]),
    .f(al_3bd314e4[64]),
    .o(al_2d07102b));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_e0588beb (
    .a(al_1634b160),
    .b(al_2d07102b),
    .c(al_3bd314e4[48]),
    .d(al_3bd314e4[49]),
    .e(al_3bd314e4[50]),
    .f(al_3bd314e4[53]),
    .o(al_3b0f07fc));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_29f34f26 (
    .a(al_3bd314e4[67]),
    .b(al_3bd314e4[68]),
    .c(al_3bd314e4[71]),
    .d(al_3bd314e4[72]),
    .e(al_3bd314e4[74]),
    .f(al_3bd314e4[77]),
    .o(al_45fda30c));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_f3198c80 (
    .a(al_3bd314e4[54]),
    .b(al_3bd314e4[57]),
    .c(al_3bd314e4[59]),
    .d(al_3bd314e4[60]),
    .e(al_3bd314e4[62]),
    .f(al_3bd314e4[65]),
    .o(al_ca8a5a31));
  AL_MAP_LUT6 #(
    .EQN("(F*~(B*A*(D@(~E*C))))"),
    .INIT(64'h77fff77f00000000))
    al_5dd7d412 (
    .a(al_3b0f07fc),
    .b(al_fd5ea84d),
    .c(al_3bd314e4[46]),
    .d(al_3bd314e4[47]),
    .e(al_83a08f3f[46]),
    .f(al_83a08f3f[47]),
    .o(al_89f2771a[47]));
  AL_DFF_X al_7c011a17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[0]));
  AL_DFF_X al_6d24de7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[9]));
  AL_DFF_X al_7a7660f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[10]));
  AL_DFF_X al_ecadcd9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[11]));
  AL_DFF_X al_f0c1c074 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[12]));
  AL_DFF_X al_a383f515 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[13]));
  AL_DFF_X al_4fd5f6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[14]));
  AL_DFF_X al_908b148d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[15]));
  AL_DFF_X al_a4edd3df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[16]));
  AL_DFF_X al_b2a6849 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[17]));
  AL_DFF_X al_fc3fe39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[18]));
  AL_DFF_X al_378853ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[1]));
  AL_DFF_X al_5dcaf2f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[19]));
  AL_DFF_X al_d624001a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[20]));
  AL_DFF_X al_5f99a6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[21]));
  AL_DFF_X al_14d76e1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[22]));
  AL_DFF_X al_44b5be7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[23]));
  AL_DFF_X al_99ac20b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[24]));
  AL_DFF_X al_968115cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[25]));
  AL_DFF_X al_826adc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[26]));
  AL_DFF_X al_4c82815 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[27]));
  AL_DFF_X al_f3e6bfb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[28]));
  AL_DFF_X al_a3af72d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[2]));
  AL_DFF_X al_b0bd650c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[29]));
  AL_DFF_X al_a29aa60e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[30]));
  AL_DFF_X al_a56ef06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[31]));
  AL_DFF_X al_eed2d6b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[32]));
  AL_DFF_X al_a0166c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[33]));
  AL_DFF_X al_e7c8ec67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[34]));
  AL_DFF_X al_8bdf8403 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[35]));
  AL_DFF_X al_5dd504c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[36]));
  AL_DFF_X al_d419daf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[37]));
  AL_DFF_X al_3328afda (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[38]));
  AL_DFF_X al_2e1eec11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[3]));
  AL_DFF_X al_4a4d438f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[39]));
  AL_DFF_X al_4d7e532d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[40]));
  AL_DFF_X al_b85ad1e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[41]));
  AL_DFF_X al_672267d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[42]));
  AL_DFF_X al_1df9fdc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[43]));
  AL_DFF_X al_6ac623e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[44]));
  AL_DFF_X al_f4a37ecf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[45]));
  AL_DFF_X al_3a0bb276 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_89f2771a[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[46]));
  AL_DFF_X al_b7d2da4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_89f2771a[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[47]));
  AL_DFF_X al_f530f996 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[4]));
  AL_DFF_X al_b0b60ff2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[5]));
  AL_DFF_X al_eecf6af9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[6]));
  AL_DFF_X al_2dcfb993 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[7]));
  AL_DFF_X al_f7e89a06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_83a08f3f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3d0cfeb4[8]));
  AL_DFF_X al_804e714f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ff28a985),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b54c1014[0]));
  AL_DFF_X al_70c9a5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_33c3313d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b54c1014[1]));
  AL_DFF_X al_ed156b68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1c8da1e8[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_acb3303d[0]));
  AL_DFF_X al_b83acd25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[26]));
  AL_DFF_X al_f2eef9e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[27]));
  AL_DFF_X al_69514422 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[28]));
  AL_DFF_X al_61c2d370 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[29]));
  AL_DFF_X al_4c9c3c0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[30]));
  AL_DFF_X al_e81551f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[31]));
  AL_DFF_X al_46173d5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[32]));
  AL_DFF_X al_4651f9c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[33]));
  AL_DFF_X al_93bf617f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[34]));
  AL_DFF_X al_34685dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[35]));
  AL_DFF_X al_ca2def8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[36]));
  AL_DFF_X al_20b84caa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[37]));
  AL_DFF_X al_2b44202c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[38]));
  AL_DFF_X al_884bdcb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[39]));
  AL_DFF_X al_5a127bfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[40]));
  AL_DFF_X al_66d93e0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[41]));
  AL_DFF_X al_b229951 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[42]));
  AL_DFF_X al_d0c2663 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[43]));
  AL_DFF_X al_58b77fa0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[44]));
  AL_DFF_X al_d13a58f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[45]));
  AL_DFF_X al_8dcec468 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[46]));
  AL_DFF_X al_38e3f590 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[47]));
  AL_DFF_X al_8e4a4f9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[48]));
  AL_DFF_X al_a4089859 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[49]));
  AL_DFF_X al_6f40b148 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[50]));
  AL_DFF_X al_d68beb89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[51]));
  AL_DFF_X al_b3944ddb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[52]));
  AL_DFF_X al_f920488f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[53]));
  AL_DFF_X al_6e64bc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[54]));
  AL_DFF_X al_96ca3016 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[55]));
  AL_DFF_X al_c296992c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[56]));
  AL_DFF_X al_19649ff2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e803eabe[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_753f5f88[57]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_b085a86b (
    .a(1'b0),
    .o({al_b8462556,open_n62}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cf8cc49e (
    .a(al_80a0f09e[27]),
    .b(al_e803eabe[27]),
    .c(al_b8462556),
    .o({al_54775a2b,al_b2ee1d57[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40bb9513 (
    .a(al_80a0f09e[28]),
    .b(al_e803eabe[28]),
    .c(al_54775a2b),
    .o({al_39d57d97,al_b2ee1d57[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6531fd23 (
    .a(al_80a0f09e[29]),
    .b(al_e803eabe[29]),
    .c(al_39d57d97),
    .o({al_e98f3c34,al_b2ee1d57[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6c13b7f2 (
    .a(al_80a0f09e[30]),
    .b(al_e803eabe[30]),
    .c(al_e98f3c34),
    .o({al_5761f230,al_b2ee1d57[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2e8683e3 (
    .a(al_80a0f09e[31]),
    .b(al_e803eabe[31]),
    .c(al_5761f230),
    .o({al_2283cfcc,al_b2ee1d57[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_43a110a4 (
    .a(al_80a0f09e[32]),
    .b(al_e803eabe[32]),
    .c(al_2283cfcc),
    .o({al_5d7328e8,al_b2ee1d57[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c879bab (
    .a(al_80a0f09e[33]),
    .b(al_e803eabe[33]),
    .c(al_5d7328e8),
    .o({al_93496304,al_b2ee1d57[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2917a840 (
    .a(al_80a0f09e[34]),
    .b(al_e803eabe[34]),
    .c(al_93496304),
    .o({al_abc34969,al_b2ee1d57[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_28cf777d (
    .a(al_80a0f09e[35]),
    .b(al_e803eabe[35]),
    .c(al_abc34969),
    .o({al_90929116,al_b2ee1d57[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_33a563e (
    .a(al_80a0f09e[36]),
    .b(al_e803eabe[36]),
    .c(al_90929116),
    .o({al_2da51efc,al_b2ee1d57[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68b0f6e (
    .a(al_80a0f09e[37]),
    .b(al_e803eabe[37]),
    .c(al_2da51efc),
    .o({al_c89089ad,al_b2ee1d57[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ded6dc50 (
    .a(al_80a0f09e[38]),
    .b(al_e803eabe[38]),
    .c(al_c89089ad),
    .o({al_e37f1d18,al_b2ee1d57[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f780a6e5 (
    .a(al_80a0f09e[39]),
    .b(al_e803eabe[39]),
    .c(al_e37f1d18),
    .o({al_77a0ba2a,al_b2ee1d57[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dee2e250 (
    .a(al_80a0f09e[40]),
    .b(al_e803eabe[40]),
    .c(al_77a0ba2a),
    .o({al_c1b434db,al_b2ee1d57[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1056452c (
    .a(al_80a0f09e[41]),
    .b(al_e803eabe[41]),
    .c(al_c1b434db),
    .o({al_5622df9b,al_b2ee1d57[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5b7f004b (
    .a(al_80a0f09e[42]),
    .b(al_e803eabe[42]),
    .c(al_5622df9b),
    .o({al_e3ce0c99,al_b2ee1d57[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cdfa7dbd (
    .a(al_80a0f09e[43]),
    .b(al_e803eabe[43]),
    .c(al_e3ce0c99),
    .o({al_7a39fd90,al_b2ee1d57[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_50e9f109 (
    .a(al_80a0f09e[44]),
    .b(al_e803eabe[44]),
    .c(al_7a39fd90),
    .o({al_290a897c,al_b2ee1d57[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1fe35401 (
    .a(al_80a0f09e[45]),
    .b(al_e803eabe[45]),
    .c(al_290a897c),
    .o({al_39495ba2,al_b2ee1d57[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4d74d3d0 (
    .a(al_80a0f09e[46]),
    .b(al_e803eabe[46]),
    .c(al_39495ba2),
    .o({al_ff8767e1,al_b2ee1d57[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc4264d9 (
    .a(al_80a0f09e[47]),
    .b(al_e803eabe[47]),
    .c(al_ff8767e1),
    .o({al_edbcd561,al_b2ee1d57[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2c291e17 (
    .c(al_edbcd561),
    .o({open_n65,al_b2ee1d57[21]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_462139c4 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[27]),
    .c(al_b2ee1d57[0]),
    .o(al_cdad9264[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9c0350ac (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[28]),
    .c(al_b2ee1d57[1]),
    .o(al_cdad9264[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_add5fc3f (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[29]),
    .c(al_b2ee1d57[2]),
    .o(al_cdad9264[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8e94977e (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[30]),
    .c(al_b2ee1d57[3]),
    .o(al_cdad9264[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_58f6f719 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[31]),
    .c(al_b2ee1d57[4]),
    .o(al_cdad9264[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a17690d3 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[32]),
    .c(al_b2ee1d57[5]),
    .o(al_cdad9264[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e34a9270 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[33]),
    .c(al_b2ee1d57[6]),
    .o(al_cdad9264[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f0ec968e (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[34]),
    .c(al_b2ee1d57[7]),
    .o(al_cdad9264[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2bfaed3d (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[35]),
    .c(al_b2ee1d57[8]),
    .o(al_cdad9264[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b226c66 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[36]),
    .c(al_b2ee1d57[9]),
    .o(al_cdad9264[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7d3865c0 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[37]),
    .c(al_b2ee1d57[10]),
    .o(al_cdad9264[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ebbc4ade (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[38]),
    .c(al_b2ee1d57[11]),
    .o(al_cdad9264[38]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_4d597a5d (
    .a(al_e803eabe[54]),
    .b(al_e803eabe[55]),
    .c(al_e803eabe[56]),
    .d(al_e803eabe[57]),
    .e(al_e803eabe[58]),
    .f(al_b2ee1d57[21]),
    .o(al_b68658c6));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_d063b6cf (
    .a(al_e803eabe[48]),
    .b(al_e803eabe[49]),
    .c(al_e803eabe[50]),
    .d(al_e803eabe[51]),
    .e(al_e803eabe[52]),
    .f(al_e803eabe[53]),
    .o(al_7bc5cf46));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_b82f2823 (
    .a(al_b68658c6),
    .b(al_7bc5cf46),
    .o(al_c9c0b8e5));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_235205ed (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[39]),
    .c(al_b2ee1d57[12]),
    .o(al_cdad9264[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ba6b069f (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[40]),
    .c(al_b2ee1d57[13]),
    .o(al_cdad9264[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_34fbf8b7 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[41]),
    .c(al_b2ee1d57[14]),
    .o(al_cdad9264[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2a42789b (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[42]),
    .c(al_b2ee1d57[15]),
    .o(al_cdad9264[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9ac2675a (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[43]),
    .c(al_b2ee1d57[16]),
    .o(al_cdad9264[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_49c440b8 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[44]),
    .c(al_b2ee1d57[17]),
    .o(al_cdad9264[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e2595a22 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[45]),
    .c(al_b2ee1d57[18]),
    .o(al_cdad9264[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_da5939bf (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[46]),
    .c(al_b2ee1d57[19]),
    .o(al_cdad9264[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_427a3d53 (
    .a(al_c9c0b8e5),
    .b(al_80a0f09e[47]),
    .c(al_b2ee1d57[20]),
    .o(al_cdad9264[47]));
  AL_DFF_X al_5320058e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[0]));
  AL_DFF_X al_81e0bd9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[9]));
  AL_DFF_X al_7dc149fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[10]));
  AL_DFF_X al_979295cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[11]));
  AL_DFF_X al_3e9b0f40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[12]));
  AL_DFF_X al_3e16e4c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[13]));
  AL_DFF_X al_6b0b9152 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[14]));
  AL_DFF_X al_2f0d228b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[15]));
  AL_DFF_X al_36f7a2d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[16]));
  AL_DFF_X al_b9b0885 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[17]));
  AL_DFF_X al_347d9dfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[18]));
  AL_DFF_X al_b6439028 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[1]));
  AL_DFF_X al_5422cb0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[19]));
  AL_DFF_X al_f29e907d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[20]));
  AL_DFF_X al_be4a1174 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[21]));
  AL_DFF_X al_77d5e301 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[22]));
  AL_DFF_X al_73ecd4d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[23]));
  AL_DFF_X al_afaee291 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[24]));
  AL_DFF_X al_f643ef18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[25]));
  AL_DFF_X al_47ac5a9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[26]));
  AL_DFF_X al_d9d77a38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[27]));
  AL_DFF_X al_55d89ae4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[28]));
  AL_DFF_X al_69b43bd6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[2]));
  AL_DFF_X al_4fdc9972 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[29]));
  AL_DFF_X al_7c0b70e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[30]));
  AL_DFF_X al_c7cc8d98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[31]));
  AL_DFF_X al_9e32cb37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[32]));
  AL_DFF_X al_e47b10cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[33]));
  AL_DFF_X al_7b08f9c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[34]));
  AL_DFF_X al_5eccc061 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[35]));
  AL_DFF_X al_5241b11f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[36]));
  AL_DFF_X al_d9fe995a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[37]));
  AL_DFF_X al_e6e00f6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[38]));
  AL_DFF_X al_df9af576 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[3]));
  AL_DFF_X al_eb4df30e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[39]));
  AL_DFF_X al_35858a73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[40]));
  AL_DFF_X al_8b8714cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[41]));
  AL_DFF_X al_b4a1a8ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[42]));
  AL_DFF_X al_df62f9fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[43]));
  AL_DFF_X al_d8bb1d4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[44]));
  AL_DFF_X al_4fff7b2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[45]));
  AL_DFF_X al_b20e6a5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[46]));
  AL_DFF_X al_b38c36ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cdad9264[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[47]));
  AL_DFF_X al_2efc7d3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[4]));
  AL_DFF_X al_650c703d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[5]));
  AL_DFF_X al_d151ad0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[6]));
  AL_DFF_X al_98779bba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[7]));
  AL_DFF_X al_171537c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_80a0f09e[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_98494645[8]));
  AL_DFF_X al_87ec2fb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c9c0b8e5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[0]));
  AL_DFF_X al_1c8d6578 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[9]));
  AL_DFF_X al_35d6e646 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[10]));
  AL_DFF_X al_ed1867b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[11]));
  AL_DFF_X al_600c496d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[12]));
  AL_DFF_X al_a8f36d24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[13]));
  AL_DFF_X al_9fb96996 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[14]));
  AL_DFF_X al_1ec0b676 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[15]));
  AL_DFF_X al_1157657d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[16]));
  AL_DFF_X al_962c0f8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[17]));
  AL_DFF_X al_36fbe55d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[18]));
  AL_DFF_X al_c57460f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[1]));
  AL_DFF_X al_49070b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[19]));
  AL_DFF_X al_1e034fc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[20]));
  AL_DFF_X al_53c6b5f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[2]));
  AL_DFF_X al_edc3444b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[3]));
  AL_DFF_X al_ad6e8ade (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[4]));
  AL_DFF_X al_e59d91d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[5]));
  AL_DFF_X al_ce2609bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[6]));
  AL_DFF_X al_54080a60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[7]));
  AL_DFF_X al_9c497eec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bd7f7f17[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_be8c4478[8]));
  AL_DFF_X al_88b2e307 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_acb3303d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_14a1a59a[0]));
  AL_DFF_X al_c05a6b81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[25]));
  AL_DFF_X al_ba406f32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[26]));
  AL_DFF_X al_a4d4b5a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[27]));
  AL_DFF_X al_c289942a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[28]));
  AL_DFF_X al_9ea39029 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[29]));
  AL_DFF_X al_af446fbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[30]));
  AL_DFF_X al_3c347408 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[31]));
  AL_DFF_X al_719d11a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[32]));
  AL_DFF_X al_13a039e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[33]));
  AL_DFF_X al_325f3245 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[34]));
  AL_DFF_X al_df3e3bd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[35]));
  AL_DFF_X al_123fa5dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[36]));
  AL_DFF_X al_431854c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[37]));
  AL_DFF_X al_6a9600a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[38]));
  AL_DFF_X al_efc43c06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[39]));
  AL_DFF_X al_1712b0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[40]));
  AL_DFF_X al_458cd162 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[41]));
  AL_DFF_X al_36a1759a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[42]));
  AL_DFF_X al_116bef1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[43]));
  AL_DFF_X al_5d2fd705 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[44]));
  AL_DFF_X al_6d692414 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[45]));
  AL_DFF_X al_2d4d3db9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[46]));
  AL_DFF_X al_7e4abe78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[47]));
  AL_DFF_X al_d93f5dcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[48]));
  AL_DFF_X al_7dc1f21e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[49]));
  AL_DFF_X al_320ee700 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[50]));
  AL_DFF_X al_b4130e4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[51]));
  AL_DFF_X al_f9282669 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[52]));
  AL_DFF_X al_e8500e88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[53]));
  AL_DFF_X al_1b3ff000 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[54]));
  AL_DFF_X al_236ce89a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[55]));
  AL_DFF_X al_16058afc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_753f5f88[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_35594bd9[56]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_6d758be1 (
    .a(1'b0),
    .o({al_ddf57730,open_n68}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c78ac8c3 (
    .a(al_98494645[26]),
    .b(al_753f5f88[26]),
    .c(al_ddf57730),
    .o({al_bcf04c60,al_3e64f540[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_58dd1907 (
    .a(al_98494645[27]),
    .b(al_753f5f88[27]),
    .c(al_bcf04c60),
    .o({al_76e6b917,al_3e64f540[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dfa782de (
    .a(al_98494645[28]),
    .b(al_753f5f88[28]),
    .c(al_76e6b917),
    .o({al_f66e0990,al_3e64f540[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a12bb745 (
    .a(al_98494645[29]),
    .b(al_753f5f88[29]),
    .c(al_f66e0990),
    .o({al_c0b6cd6e,al_3e64f540[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a0885ec5 (
    .a(al_98494645[30]),
    .b(al_753f5f88[30]),
    .c(al_c0b6cd6e),
    .o({al_5507d757,al_3e64f540[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f8bda533 (
    .a(al_98494645[31]),
    .b(al_753f5f88[31]),
    .c(al_5507d757),
    .o({al_216ce40,al_3e64f540[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4c6baf49 (
    .a(al_98494645[32]),
    .b(al_753f5f88[32]),
    .c(al_216ce40),
    .o({al_66aff298,al_3e64f540[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ec721979 (
    .a(al_98494645[33]),
    .b(al_753f5f88[33]),
    .c(al_66aff298),
    .o({al_cdeed011,al_3e64f540[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ad96c833 (
    .a(al_98494645[34]),
    .b(al_753f5f88[34]),
    .c(al_cdeed011),
    .o({al_d2fa64e6,al_3e64f540[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_36c06626 (
    .a(al_98494645[35]),
    .b(al_753f5f88[35]),
    .c(al_d2fa64e6),
    .o({al_e0707d5b,al_3e64f540[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_79fe47b8 (
    .a(al_98494645[36]),
    .b(al_753f5f88[36]),
    .c(al_e0707d5b),
    .o({al_b9091bb4,al_3e64f540[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67f00340 (
    .a(al_98494645[37]),
    .b(al_753f5f88[37]),
    .c(al_b9091bb4),
    .o({al_cafa3568,al_3e64f540[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6cedabdb (
    .a(al_98494645[38]),
    .b(al_753f5f88[38]),
    .c(al_cafa3568),
    .o({al_177f9d69,al_3e64f540[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_382e81bd (
    .a(al_98494645[39]),
    .b(al_753f5f88[39]),
    .c(al_177f9d69),
    .o({al_8d529875,al_3e64f540[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5b66c624 (
    .a(al_98494645[40]),
    .b(al_753f5f88[40]),
    .c(al_8d529875),
    .o({al_663d37b6,al_3e64f540[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bd56bc0 (
    .a(al_98494645[41]),
    .b(al_753f5f88[41]),
    .c(al_663d37b6),
    .o({al_bd5caa9f,al_3e64f540[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b30895d (
    .a(al_98494645[42]),
    .b(al_753f5f88[42]),
    .c(al_bd5caa9f),
    .o({al_95b12900,al_3e64f540[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_82c9ab03 (
    .a(al_98494645[43]),
    .b(al_753f5f88[43]),
    .c(al_95b12900),
    .o({al_a9d8f8,al_3e64f540[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e29bec0b (
    .a(al_98494645[44]),
    .b(al_753f5f88[44]),
    .c(al_a9d8f8),
    .o({al_3459937f,al_3e64f540[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b28007b (
    .a(al_98494645[45]),
    .b(al_753f5f88[45]),
    .c(al_3459937f),
    .o({al_b062dbda,al_3e64f540[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_689c8fae (
    .a(al_98494645[46]),
    .b(al_753f5f88[46]),
    .c(al_b062dbda),
    .o({al_ab1c35b3,al_3e64f540[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b7429878 (
    .a(al_98494645[47]),
    .b(al_753f5f88[47]),
    .c(al_ab1c35b3),
    .o({al_41371141,al_3e64f540[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67de1a93 (
    .c(al_41371141),
    .o({open_n71,al_3e64f540[22]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_18f302d2 (
    .a(al_8f25dca0),
    .b(al_98494645[26]),
    .c(al_3e64f540[0]),
    .o(al_f7ed724c[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c538154a (
    .a(al_8f25dca0),
    .b(al_98494645[27]),
    .c(al_3e64f540[1]),
    .o(al_f7ed724c[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e08f281b (
    .a(al_8f25dca0),
    .b(al_98494645[28]),
    .c(al_3e64f540[2]),
    .o(al_f7ed724c[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_99561eae (
    .a(al_8f25dca0),
    .b(al_98494645[29]),
    .c(al_3e64f540[3]),
    .o(al_f7ed724c[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_369dde19 (
    .a(al_8f25dca0),
    .b(al_98494645[30]),
    .c(al_3e64f540[4]),
    .o(al_f7ed724c[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2e402e97 (
    .a(al_8f25dca0),
    .b(al_98494645[31]),
    .c(al_3e64f540[5]),
    .o(al_f7ed724c[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_df41b7d4 (
    .a(al_8f25dca0),
    .b(al_98494645[32]),
    .c(al_3e64f540[6]),
    .o(al_f7ed724c[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cb82d410 (
    .a(al_8f25dca0),
    .b(al_98494645[33]),
    .c(al_3e64f540[7]),
    .o(al_f7ed724c[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e66781f0 (
    .a(al_8f25dca0),
    .b(al_98494645[34]),
    .c(al_3e64f540[8]),
    .o(al_f7ed724c[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e4560ea1 (
    .a(al_8f25dca0),
    .b(al_98494645[35]),
    .c(al_3e64f540[9]),
    .o(al_f7ed724c[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_40401160 (
    .a(al_8f25dca0),
    .b(al_98494645[36]),
    .c(al_3e64f540[10]),
    .o(al_f7ed724c[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_598a9821 (
    .a(al_8f25dca0),
    .b(al_98494645[37]),
    .c(al_3e64f540[11]),
    .o(al_f7ed724c[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_82fc2728 (
    .a(al_8f25dca0),
    .b(al_98494645[38]),
    .c(al_3e64f540[12]),
    .o(al_f7ed724c[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_20a8f0dc (
    .a(al_8f25dca0),
    .b(al_98494645[39]),
    .c(al_3e64f540[13]),
    .o(al_f7ed724c[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_51a28816 (
    .a(al_8f25dca0),
    .b(al_98494645[40]),
    .c(al_3e64f540[14]),
    .o(al_f7ed724c[40]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_de834657 (
    .a(al_753f5f88[52]),
    .b(al_753f5f88[53]),
    .c(al_753f5f88[54]),
    .d(al_753f5f88[55]),
    .e(al_753f5f88[56]),
    .f(al_753f5f88[57]),
    .o(al_a7492340));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*A)"),
    .INIT(64'h0000000000000002))
    al_cfcf42c1 (
    .a(al_a7492340),
    .b(al_753f5f88[48]),
    .c(al_753f5f88[49]),
    .d(al_753f5f88[50]),
    .e(al_753f5f88[51]),
    .f(al_3e64f540[22]),
    .o(al_8f25dca0));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_73cd6c47 (
    .a(al_8f25dca0),
    .b(al_98494645[41]),
    .c(al_3e64f540[15]),
    .o(al_f7ed724c[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_de126eba (
    .a(al_8f25dca0),
    .b(al_98494645[42]),
    .c(al_3e64f540[16]),
    .o(al_f7ed724c[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8d864ae7 (
    .a(al_8f25dca0),
    .b(al_98494645[43]),
    .c(al_3e64f540[17]),
    .o(al_f7ed724c[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e548b7f8 (
    .a(al_8f25dca0),
    .b(al_98494645[44]),
    .c(al_3e64f540[18]),
    .o(al_f7ed724c[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8e72051e (
    .a(al_8f25dca0),
    .b(al_98494645[45]),
    .c(al_3e64f540[19]),
    .o(al_f7ed724c[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_81c51432 (
    .a(al_8f25dca0),
    .b(al_98494645[46]),
    .c(al_3e64f540[20]),
    .o(al_f7ed724c[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7b8c2610 (
    .a(al_8f25dca0),
    .b(al_98494645[47]),
    .c(al_3e64f540[21]),
    .o(al_f7ed724c[47]));
  AL_DFF_X al_bb3f5483 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[0]));
  AL_DFF_X al_c8f15ee8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[9]));
  AL_DFF_X al_a7fddae4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[10]));
  AL_DFF_X al_6c911d7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[11]));
  AL_DFF_X al_983b8d7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[12]));
  AL_DFF_X al_4aa9eff0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[13]));
  AL_DFF_X al_f6707563 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[14]));
  AL_DFF_X al_d83bb58e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[15]));
  AL_DFF_X al_ce23af80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[16]));
  AL_DFF_X al_6eb8b053 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[17]));
  AL_DFF_X al_37eda87c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[18]));
  AL_DFF_X al_9d43c75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[1]));
  AL_DFF_X al_d15ad720 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[19]));
  AL_DFF_X al_de54bf66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[20]));
  AL_DFF_X al_b79f1af5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[21]));
  AL_DFF_X al_3350f0d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[22]));
  AL_DFF_X al_f380a039 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[23]));
  AL_DFF_X al_1d7792d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[24]));
  AL_DFF_X al_5d6904fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[25]));
  AL_DFF_X al_d498611b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[26]));
  AL_DFF_X al_25ce006b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[27]));
  AL_DFF_X al_f5740c40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[28]));
  AL_DFF_X al_47f9b70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[2]));
  AL_DFF_X al_64c7122f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[29]));
  AL_DFF_X al_5c7ae4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[30]));
  AL_DFF_X al_8d97b054 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[31]));
  AL_DFF_X al_fda37d80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[32]));
  AL_DFF_X al_b4176e97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[33]));
  AL_DFF_X al_c1b411c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[34]));
  AL_DFF_X al_801e8e9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[35]));
  AL_DFF_X al_a6ac9ed9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[36]));
  AL_DFF_X al_d671d436 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[37]));
  AL_DFF_X al_90db964d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[38]));
  AL_DFF_X al_e9adc848 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[3]));
  AL_DFF_X al_d0842f97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[39]));
  AL_DFF_X al_26b6d7ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[40]));
  AL_DFF_X al_d8a37af5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[41]));
  AL_DFF_X al_65a64e74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[42]));
  AL_DFF_X al_3a620b45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[43]));
  AL_DFF_X al_dce4fa5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[44]));
  AL_DFF_X al_6e15a454 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[45]));
  AL_DFF_X al_15248ded (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[46]));
  AL_DFF_X al_b90e5663 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7ed724c[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[47]));
  AL_DFF_X al_b69591be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[4]));
  AL_DFF_X al_87b5e23d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[5]));
  AL_DFF_X al_2620849d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[6]));
  AL_DFF_X al_d9cd4be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[7]));
  AL_DFF_X al_456cf9ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_98494645[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bf34d64d[8]));
  AL_DFF_X al_a7b45e7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8f25dca0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[0]));
  AL_DFF_X al_ea703c1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[9]));
  AL_DFF_X al_b13fefc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[10]));
  AL_DFF_X al_3f838dae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[11]));
  AL_DFF_X al_fede49ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[12]));
  AL_DFF_X al_698da4ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[13]));
  AL_DFF_X al_7190ccff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[14]));
  AL_DFF_X al_564dd794 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[15]));
  AL_DFF_X al_5dd0e62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[16]));
  AL_DFF_X al_6b743b95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[17]));
  AL_DFF_X al_31016250 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[18]));
  AL_DFF_X al_8a368b0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[1]));
  AL_DFF_X al_5239e539 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[19]));
  AL_DFF_X al_805068dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[20]));
  AL_DFF_X al_5bac1c57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[21]));
  AL_DFF_X al_375954b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[2]));
  AL_DFF_X al_52580f39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[3]));
  AL_DFF_X al_da99564e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[4]));
  AL_DFF_X al_4af5ce86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[5]));
  AL_DFF_X al_905182c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[6]));
  AL_DFF_X al_81d7a9a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[7]));
  AL_DFF_X al_f2e61415 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be8c4478[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f1d740ba[8]));
  AL_DFF_X al_5f284f64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14a1a59a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_21143207[0]));
  AL_DFF_X al_b2a5247f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[24]));
  AL_DFF_X al_a8aed8f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[25]));
  AL_DFF_X al_fbd0ed2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[26]));
  AL_DFF_X al_e167fea3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[27]));
  AL_DFF_X al_5a5577ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[28]));
  AL_DFF_X al_8616d62d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[29]));
  AL_DFF_X al_50e49a5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[30]));
  AL_DFF_X al_e99db947 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[31]));
  AL_DFF_X al_ca109159 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[32]));
  AL_DFF_X al_929daa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[33]));
  AL_DFF_X al_1d410e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[34]));
  AL_DFF_X al_4eb3563e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[35]));
  AL_DFF_X al_85fc8f6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[36]));
  AL_DFF_X al_75f6df94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[37]));
  AL_DFF_X al_6d54c6f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[38]));
  AL_DFF_X al_39c1280c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[39]));
  AL_DFF_X al_a0f84fd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[40]));
  AL_DFF_X al_4e6d1b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[41]));
  AL_DFF_X al_f15fe143 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[42]));
  AL_DFF_X al_8d2d2880 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[43]));
  AL_DFF_X al_89c0be39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[44]));
  AL_DFF_X al_98d35a48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[45]));
  AL_DFF_X al_5e8a29c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[46]));
  AL_DFF_X al_d297c1f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[47]));
  AL_DFF_X al_97cbcadb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[48]));
  AL_DFF_X al_1771ca1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[49]));
  AL_DFF_X al_a1868725 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[50]));
  AL_DFF_X al_f9717522 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[51]));
  AL_DFF_X al_3c679c1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[52]));
  AL_DFF_X al_3fec7673 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[53]));
  AL_DFF_X al_840497bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[54]));
  AL_DFF_X al_1e4035de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_35594bd9[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2bb4ec4[55]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_fc2be15c (
    .a(1'b0),
    .o({al_b27b3769,open_n74}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_af1531a2 (
    .a(al_bf34d64d[25]),
    .b(al_35594bd9[25]),
    .c(al_b27b3769),
    .o({al_a8fb6998,al_365f90b4[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_19239a5b (
    .a(al_bf34d64d[26]),
    .b(al_35594bd9[26]),
    .c(al_a8fb6998),
    .o({al_18a0a383,al_365f90b4[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ad607d9f (
    .a(al_bf34d64d[27]),
    .b(al_35594bd9[27]),
    .c(al_18a0a383),
    .o({al_2f3a1692,al_365f90b4[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f1035696 (
    .a(al_bf34d64d[28]),
    .b(al_35594bd9[28]),
    .c(al_2f3a1692),
    .o({al_d4bc7f3e,al_365f90b4[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b908b684 (
    .a(al_bf34d64d[29]),
    .b(al_35594bd9[29]),
    .c(al_d4bc7f3e),
    .o({al_72d62b1c,al_365f90b4[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_839478a1 (
    .a(al_bf34d64d[30]),
    .b(al_35594bd9[30]),
    .c(al_72d62b1c),
    .o({al_4e56a0da,al_365f90b4[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_444ba3b9 (
    .a(al_bf34d64d[31]),
    .b(al_35594bd9[31]),
    .c(al_4e56a0da),
    .o({al_1240f9a6,al_365f90b4[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4e7271bc (
    .a(al_bf34d64d[32]),
    .b(al_35594bd9[32]),
    .c(al_1240f9a6),
    .o({al_2ec3de14,al_365f90b4[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a7de056e (
    .a(al_bf34d64d[33]),
    .b(al_35594bd9[33]),
    .c(al_2ec3de14),
    .o({al_b48c402a,al_365f90b4[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee011bb9 (
    .a(al_bf34d64d[34]),
    .b(al_35594bd9[34]),
    .c(al_b48c402a),
    .o({al_63f814e,al_365f90b4[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fa7dcc79 (
    .a(al_bf34d64d[35]),
    .b(al_35594bd9[35]),
    .c(al_63f814e),
    .o({al_3c4a2199,al_365f90b4[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2c1c2419 (
    .a(al_bf34d64d[36]),
    .b(al_35594bd9[36]),
    .c(al_3c4a2199),
    .o({al_f832136c,al_365f90b4[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_97d166cd (
    .a(al_bf34d64d[37]),
    .b(al_35594bd9[37]),
    .c(al_f832136c),
    .o({al_934e501,al_365f90b4[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a9125f03 (
    .a(al_bf34d64d[38]),
    .b(al_35594bd9[38]),
    .c(al_934e501),
    .o({al_d460c819,al_365f90b4[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d612153b (
    .a(al_bf34d64d[39]),
    .b(al_35594bd9[39]),
    .c(al_d460c819),
    .o({al_88e1bda3,al_365f90b4[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b935815 (
    .a(al_bf34d64d[40]),
    .b(al_35594bd9[40]),
    .c(al_88e1bda3),
    .o({al_1821d93d,al_365f90b4[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_89b9e811 (
    .a(al_bf34d64d[41]),
    .b(al_35594bd9[41]),
    .c(al_1821d93d),
    .o({al_b4ee9e86,al_365f90b4[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dbfb13db (
    .a(al_bf34d64d[42]),
    .b(al_35594bd9[42]),
    .c(al_b4ee9e86),
    .o({al_9828f0b3,al_365f90b4[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c90a3347 (
    .a(al_bf34d64d[43]),
    .b(al_35594bd9[43]),
    .c(al_9828f0b3),
    .o({al_3f6c8445,al_365f90b4[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_893284b6 (
    .a(al_bf34d64d[44]),
    .b(al_35594bd9[44]),
    .c(al_3f6c8445),
    .o({al_28e359b1,al_365f90b4[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ae6c4b0 (
    .a(al_bf34d64d[45]),
    .b(al_35594bd9[45]),
    .c(al_28e359b1),
    .o({al_4b337999,al_365f90b4[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_37a9453a (
    .a(al_bf34d64d[46]),
    .b(al_35594bd9[46]),
    .c(al_4b337999),
    .o({al_92297df8,al_365f90b4[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_357322b7 (
    .a(al_bf34d64d[47]),
    .b(al_35594bd9[47]),
    .c(al_92297df8),
    .o({al_7dcd3618,al_365f90b4[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c12e03b3 (
    .c(al_7dcd3618),
    .o({open_n77,al_365f90b4[23]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c8755677 (
    .a(al_274f6baa),
    .b(al_bf34d64d[25]),
    .c(al_365f90b4[0]),
    .o(al_96533024[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_15a71cc6 (
    .a(al_274f6baa),
    .b(al_bf34d64d[26]),
    .c(al_365f90b4[1]),
    .o(al_96533024[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_85d5f343 (
    .a(al_274f6baa),
    .b(al_bf34d64d[27]),
    .c(al_365f90b4[2]),
    .o(al_96533024[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dfe9fd59 (
    .a(al_274f6baa),
    .b(al_bf34d64d[28]),
    .c(al_365f90b4[3]),
    .o(al_96533024[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4f01e5bc (
    .a(al_274f6baa),
    .b(al_bf34d64d[29]),
    .c(al_365f90b4[4]),
    .o(al_96533024[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d4c47521 (
    .a(al_274f6baa),
    .b(al_bf34d64d[30]),
    .c(al_365f90b4[5]),
    .o(al_96533024[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b1a091eb (
    .a(al_274f6baa),
    .b(al_bf34d64d[31]),
    .c(al_365f90b4[6]),
    .o(al_96533024[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f30ec840 (
    .a(al_274f6baa),
    .b(al_bf34d64d[32]),
    .c(al_365f90b4[7]),
    .o(al_96533024[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2832786c (
    .a(al_274f6baa),
    .b(al_bf34d64d[33]),
    .c(al_365f90b4[8]),
    .o(al_96533024[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_90fb2bc3 (
    .a(al_274f6baa),
    .b(al_bf34d64d[34]),
    .c(al_365f90b4[9]),
    .o(al_96533024[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8625cce7 (
    .a(al_274f6baa),
    .b(al_bf34d64d[35]),
    .c(al_365f90b4[10]),
    .o(al_96533024[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_59e7bdd7 (
    .a(al_274f6baa),
    .b(al_bf34d64d[36]),
    .c(al_365f90b4[11]),
    .o(al_96533024[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2e7a287f (
    .a(al_274f6baa),
    .b(al_bf34d64d[37]),
    .c(al_365f90b4[12]),
    .o(al_96533024[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4af9a9bb (
    .a(al_274f6baa),
    .b(al_bf34d64d[38]),
    .c(al_365f90b4[13]),
    .o(al_96533024[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bab67d18 (
    .a(al_274f6baa),
    .b(al_bf34d64d[39]),
    .c(al_365f90b4[14]),
    .o(al_96533024[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8e74cbbe (
    .a(al_274f6baa),
    .b(al_bf34d64d[40]),
    .c(al_365f90b4[15]),
    .o(al_96533024[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e67163f (
    .a(al_274f6baa),
    .b(al_bf34d64d[41]),
    .c(al_365f90b4[16]),
    .o(al_96533024[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_53b7b84e (
    .a(al_274f6baa),
    .b(al_bf34d64d[42]),
    .c(al_365f90b4[17]),
    .o(al_96533024[42]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_377cce25 (
    .a(al_35594bd9[52]),
    .b(al_35594bd9[53]),
    .c(al_35594bd9[54]),
    .d(al_35594bd9[55]),
    .e(al_35594bd9[56]),
    .f(al_365f90b4[23]),
    .o(al_68deb8d6));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    al_9bda22d5 (
    .a(al_68deb8d6),
    .b(al_35594bd9[48]),
    .c(al_35594bd9[49]),
    .d(al_35594bd9[50]),
    .e(al_35594bd9[51]),
    .o(al_274f6baa));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fe63cf35 (
    .a(al_274f6baa),
    .b(al_bf34d64d[43]),
    .c(al_365f90b4[18]),
    .o(al_96533024[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_38fce98c (
    .a(al_274f6baa),
    .b(al_bf34d64d[44]),
    .c(al_365f90b4[19]),
    .o(al_96533024[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b9473c5f (
    .a(al_274f6baa),
    .b(al_bf34d64d[45]),
    .c(al_365f90b4[20]),
    .o(al_96533024[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f1011bca (
    .a(al_274f6baa),
    .b(al_bf34d64d[46]),
    .c(al_365f90b4[21]),
    .o(al_96533024[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_45b4a74b (
    .a(al_274f6baa),
    .b(al_bf34d64d[47]),
    .c(al_365f90b4[22]),
    .o(al_96533024[47]));
  AL_DFF_X al_d8052def (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[0]));
  AL_DFF_X al_f6daf26f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[9]));
  AL_DFF_X al_44a614a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[10]));
  AL_DFF_X al_55f95e93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[11]));
  AL_DFF_X al_5dfc1670 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[12]));
  AL_DFF_X al_c4ae9a74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[13]));
  AL_DFF_X al_fc4bfccc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[14]));
  AL_DFF_X al_b90baf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[15]));
  AL_DFF_X al_6acc24cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[16]));
  AL_DFF_X al_b7cf4adb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[17]));
  AL_DFF_X al_8b708de5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[18]));
  AL_DFF_X al_2b750f9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[1]));
  AL_DFF_X al_bf33a2d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[19]));
  AL_DFF_X al_913b80b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[20]));
  AL_DFF_X al_a9f7368c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[21]));
  AL_DFF_X al_942b6ce5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[22]));
  AL_DFF_X al_4fe7f524 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[23]));
  AL_DFF_X al_ba79f0a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[24]));
  AL_DFF_X al_2c6ebf10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[25]));
  AL_DFF_X al_5631130f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[26]));
  AL_DFF_X al_f9301824 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[27]));
  AL_DFF_X al_2b90b67f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[28]));
  AL_DFF_X al_6d8fc268 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[2]));
  AL_DFF_X al_dd318899 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[29]));
  AL_DFF_X al_c1571600 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[30]));
  AL_DFF_X al_9def1109 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[31]));
  AL_DFF_X al_3eb3ce4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[32]));
  AL_DFF_X al_79ef3beb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[33]));
  AL_DFF_X al_6765672 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[34]));
  AL_DFF_X al_90cd1050 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[35]));
  AL_DFF_X al_7593f9a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[36]));
  AL_DFF_X al_c98f44ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[37]));
  AL_DFF_X al_68e1c075 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[38]));
  AL_DFF_X al_205ec69c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[3]));
  AL_DFF_X al_e83acc24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[39]));
  AL_DFF_X al_8cbe24ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[40]));
  AL_DFF_X al_91ab386b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[41]));
  AL_DFF_X al_84c92c1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[42]));
  AL_DFF_X al_1aa6c4c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[43]));
  AL_DFF_X al_ca758aa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[44]));
  AL_DFF_X al_debacbbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[45]));
  AL_DFF_X al_86d9c240 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[46]));
  AL_DFF_X al_15abf01e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_96533024[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[47]));
  AL_DFF_X al_930a9639 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[4]));
  AL_DFF_X al_896f2461 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[5]));
  AL_DFF_X al_69d8e945 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[6]));
  AL_DFF_X al_7dcb3a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[7]));
  AL_DFF_X al_3b51a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bf34d64d[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f0f43754[8]));
  AL_DFF_X al_3524e5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_274f6baa),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[0]));
  AL_DFF_X al_92edde8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[9]));
  AL_DFF_X al_976eab0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[10]));
  AL_DFF_X al_ab26d617 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[11]));
  AL_DFF_X al_7bba285f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[12]));
  AL_DFF_X al_7c45a303 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[13]));
  AL_DFF_X al_a4e0d6a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[14]));
  AL_DFF_X al_f19e78da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[15]));
  AL_DFF_X al_abc7ac54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[16]));
  AL_DFF_X al_2d352fe4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[17]));
  AL_DFF_X al_4237fa9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[18]));
  AL_DFF_X al_f6303539 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[1]));
  AL_DFF_X al_812d4af7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[19]));
  AL_DFF_X al_c7402da0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[20]));
  AL_DFF_X al_d2da92a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[21]));
  AL_DFF_X al_35fcd002 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[22]));
  AL_DFF_X al_19927e4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[2]));
  AL_DFF_X al_fab6cb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[3]));
  AL_DFF_X al_e2a7c7ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[4]));
  AL_DFF_X al_b05763e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[5]));
  AL_DFF_X al_65eec0df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[6]));
  AL_DFF_X al_5e1fca8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[7]));
  AL_DFF_X al_eca117a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f1d740ba[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d3734717[8]));
  AL_DFF_X al_9979266b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_21143207[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e0dc7e9e[0]));
  AL_DFF_X al_323e68ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[23]));
  AL_DFF_X al_f7701d66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[24]));
  AL_DFF_X al_9f0b5dc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[25]));
  AL_DFF_X al_193fd2cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[26]));
  AL_DFF_X al_95271a41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[27]));
  AL_DFF_X al_8851bc0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[28]));
  AL_DFF_X al_c07cec19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[29]));
  AL_DFF_X al_eeaffa73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[30]));
  AL_DFF_X al_e55bbe3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[31]));
  AL_DFF_X al_2191dcb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[32]));
  AL_DFF_X al_707aceba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[33]));
  AL_DFF_X al_e2bc48af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[34]));
  AL_DFF_X al_387f764f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[35]));
  AL_DFF_X al_a5c9ef21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[36]));
  AL_DFF_X al_9b908156 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[37]));
  AL_DFF_X al_97db4f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[38]));
  AL_DFF_X al_5f36e75e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[39]));
  AL_DFF_X al_b5009363 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[40]));
  AL_DFF_X al_5e9ff11b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[41]));
  AL_DFF_X al_3f75c2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[42]));
  AL_DFF_X al_ab2cd9b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[43]));
  AL_DFF_X al_aa0c27ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[44]));
  AL_DFF_X al_452acfd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[45]));
  AL_DFF_X al_51b50e88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[46]));
  AL_DFF_X al_b8f8bdb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[47]));
  AL_DFF_X al_4858f68a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[48]));
  AL_DFF_X al_5a0d9df1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[49]));
  AL_DFF_X al_a27f890a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[50]));
  AL_DFF_X al_8e144b6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[51]));
  AL_DFF_X al_d4567b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[52]));
  AL_DFF_X al_799e615 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[53]));
  AL_DFF_X al_9fc4c0db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2bb4ec4[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3029c49a[54]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_253239be (
    .a(1'b0),
    .o({al_86dc2d65,open_n80}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_54b339de (
    .a(al_f0f43754[24]),
    .b(al_f2bb4ec4[24]),
    .c(al_86dc2d65),
    .o({al_f4230bb8,al_21ee8bc[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a93408b (
    .a(al_f0f43754[25]),
    .b(al_f2bb4ec4[25]),
    .c(al_f4230bb8),
    .o({al_ada1b083,al_21ee8bc[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7d0a4b60 (
    .a(al_f0f43754[26]),
    .b(al_f2bb4ec4[26]),
    .c(al_ada1b083),
    .o({al_5051b702,al_21ee8bc[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd65ddfc (
    .a(al_f0f43754[27]),
    .b(al_f2bb4ec4[27]),
    .c(al_5051b702),
    .o({al_fd100c07,al_21ee8bc[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_56ddef48 (
    .a(al_f0f43754[28]),
    .b(al_f2bb4ec4[28]),
    .c(al_fd100c07),
    .o({al_f492d664,al_21ee8bc[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1e4adae5 (
    .a(al_f0f43754[29]),
    .b(al_f2bb4ec4[29]),
    .c(al_f492d664),
    .o({al_6d3aa56f,al_21ee8bc[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc5ef7f9 (
    .a(al_f0f43754[30]),
    .b(al_f2bb4ec4[30]),
    .c(al_6d3aa56f),
    .o({al_534497b1,al_21ee8bc[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_696c4df9 (
    .a(al_f0f43754[31]),
    .b(al_f2bb4ec4[31]),
    .c(al_534497b1),
    .o({al_cb73325b,al_21ee8bc[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b29a9270 (
    .a(al_f0f43754[32]),
    .b(al_f2bb4ec4[32]),
    .c(al_cb73325b),
    .o({al_b65c9b4,al_21ee8bc[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cecd159a (
    .a(al_f0f43754[33]),
    .b(al_f2bb4ec4[33]),
    .c(al_b65c9b4),
    .o({al_178c71f6,al_21ee8bc[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_777c58f6 (
    .a(al_f0f43754[34]),
    .b(al_f2bb4ec4[34]),
    .c(al_178c71f6),
    .o({al_cbbef4f,al_21ee8bc[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_63a2c892 (
    .a(al_f0f43754[35]),
    .b(al_f2bb4ec4[35]),
    .c(al_cbbef4f),
    .o({al_9e9b738f,al_21ee8bc[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9267e288 (
    .a(al_f0f43754[36]),
    .b(al_f2bb4ec4[36]),
    .c(al_9e9b738f),
    .o({al_a076256b,al_21ee8bc[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_13389a15 (
    .a(al_f0f43754[37]),
    .b(al_f2bb4ec4[37]),
    .c(al_a076256b),
    .o({al_7930e629,al_21ee8bc[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_47728096 (
    .a(al_f0f43754[38]),
    .b(al_f2bb4ec4[38]),
    .c(al_7930e629),
    .o({al_a521f9f,al_21ee8bc[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5ef1d102 (
    .a(al_f0f43754[39]),
    .b(al_f2bb4ec4[39]),
    .c(al_a521f9f),
    .o({al_5f29b438,al_21ee8bc[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_39c0b869 (
    .a(al_f0f43754[40]),
    .b(al_f2bb4ec4[40]),
    .c(al_5f29b438),
    .o({al_3ce4b2fd,al_21ee8bc[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bd0ba43c (
    .a(al_f0f43754[41]),
    .b(al_f2bb4ec4[41]),
    .c(al_3ce4b2fd),
    .o({al_86766b99,al_21ee8bc[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6ba2c4c (
    .a(al_f0f43754[42]),
    .b(al_f2bb4ec4[42]),
    .c(al_86766b99),
    .o({al_b17e5f2d,al_21ee8bc[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_217a3a9a (
    .a(al_f0f43754[43]),
    .b(al_f2bb4ec4[43]),
    .c(al_b17e5f2d),
    .o({al_a2b56c4c,al_21ee8bc[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fe1a61c8 (
    .a(al_f0f43754[44]),
    .b(al_f2bb4ec4[44]),
    .c(al_a2b56c4c),
    .o({al_998abf81,al_21ee8bc[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_19bf4928 (
    .a(al_f0f43754[45]),
    .b(al_f2bb4ec4[45]),
    .c(al_998abf81),
    .o({al_ce61dd12,al_21ee8bc[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_526ff6eb (
    .a(al_f0f43754[46]),
    .b(al_f2bb4ec4[46]),
    .c(al_ce61dd12),
    .o({al_1ae1e567,al_21ee8bc[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6f35b9e3 (
    .a(al_f0f43754[47]),
    .b(al_f2bb4ec4[47]),
    .c(al_1ae1e567),
    .o({al_eea1c0b5,al_21ee8bc[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bb1bb8c4 (
    .c(al_eea1c0b5),
    .o({open_n83,al_21ee8bc[24]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2fbc7b03 (
    .a(al_92faecea),
    .b(al_f0f43754[24]),
    .c(al_21ee8bc[0]),
    .o(al_e60d8647[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d796eadb (
    .a(al_92faecea),
    .b(al_f0f43754[25]),
    .c(al_21ee8bc[1]),
    .o(al_e60d8647[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b4f8857c (
    .a(al_92faecea),
    .b(al_f0f43754[26]),
    .c(al_21ee8bc[2]),
    .o(al_e60d8647[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e6253bca (
    .a(al_92faecea),
    .b(al_f0f43754[27]),
    .c(al_21ee8bc[3]),
    .o(al_e60d8647[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c9732bef (
    .a(al_92faecea),
    .b(al_f0f43754[28]),
    .c(al_21ee8bc[4]),
    .o(al_e60d8647[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1491d4b7 (
    .a(al_92faecea),
    .b(al_f0f43754[29]),
    .c(al_21ee8bc[5]),
    .o(al_e60d8647[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9c82427f (
    .a(al_92faecea),
    .b(al_f0f43754[30]),
    .c(al_21ee8bc[6]),
    .o(al_e60d8647[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_47cb7671 (
    .a(al_92faecea),
    .b(al_f0f43754[31]),
    .c(al_21ee8bc[7]),
    .o(al_e60d8647[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a7cf6a44 (
    .a(al_92faecea),
    .b(al_f0f43754[32]),
    .c(al_21ee8bc[8]),
    .o(al_e60d8647[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b42b6e70 (
    .a(al_92faecea),
    .b(al_f0f43754[33]),
    .c(al_21ee8bc[9]),
    .o(al_e60d8647[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_60b076eb (
    .a(al_92faecea),
    .b(al_f0f43754[34]),
    .c(al_21ee8bc[10]),
    .o(al_e60d8647[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ba9f44e8 (
    .a(al_92faecea),
    .b(al_f0f43754[35]),
    .c(al_21ee8bc[11]),
    .o(al_e60d8647[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c3be38e1 (
    .a(al_92faecea),
    .b(al_f0f43754[36]),
    .c(al_21ee8bc[12]),
    .o(al_e60d8647[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6da340b2 (
    .a(al_92faecea),
    .b(al_f0f43754[37]),
    .c(al_21ee8bc[13]),
    .o(al_e60d8647[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b4917799 (
    .a(al_92faecea),
    .b(al_f0f43754[38]),
    .c(al_21ee8bc[14]),
    .o(al_e60d8647[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3fcf9b0d (
    .a(al_92faecea),
    .b(al_f0f43754[39]),
    .c(al_21ee8bc[15]),
    .o(al_e60d8647[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c94bd55 (
    .a(al_92faecea),
    .b(al_f0f43754[40]),
    .c(al_21ee8bc[16]),
    .o(al_e60d8647[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_18e54c80 (
    .a(al_92faecea),
    .b(al_f0f43754[41]),
    .c(al_21ee8bc[17]),
    .o(al_e60d8647[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3f1a96a (
    .a(al_92faecea),
    .b(al_f0f43754[42]),
    .c(al_21ee8bc[18]),
    .o(al_e60d8647[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_732f3f5e (
    .a(al_92faecea),
    .b(al_f0f43754[43]),
    .c(al_21ee8bc[19]),
    .o(al_e60d8647[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_395b5264 (
    .a(al_92faecea),
    .b(al_f0f43754[44]),
    .c(al_21ee8bc[20]),
    .o(al_e60d8647[44]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_274eba16 (
    .a(al_f2bb4ec4[50]),
    .b(al_f2bb4ec4[51]),
    .c(al_f2bb4ec4[52]),
    .d(al_f2bb4ec4[53]),
    .e(al_f2bb4ec4[54]),
    .f(al_f2bb4ec4[55]),
    .o(al_8d1ae89a));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    al_106d01a4 (
    .a(al_8d1ae89a),
    .b(al_f2bb4ec4[48]),
    .c(al_f2bb4ec4[49]),
    .d(al_21ee8bc[24]),
    .o(al_92faecea));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_15ce719 (
    .a(al_92faecea),
    .b(al_f0f43754[45]),
    .c(al_21ee8bc[21]),
    .o(al_e60d8647[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5e167fe (
    .a(al_92faecea),
    .b(al_f0f43754[46]),
    .c(al_21ee8bc[22]),
    .o(al_e60d8647[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_78254971 (
    .a(al_92faecea),
    .b(al_f0f43754[47]),
    .c(al_21ee8bc[23]),
    .o(al_e60d8647[47]));
  AL_DFF_X al_f4dab01f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[0]));
  AL_DFF_X al_824b1339 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[9]));
  AL_DFF_X al_a65f6058 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[10]));
  AL_DFF_X al_c51c3561 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[11]));
  AL_DFF_X al_a9d37c4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[12]));
  AL_DFF_X al_77536ad8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[13]));
  AL_DFF_X al_c9608411 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[14]));
  AL_DFF_X al_e64254f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[15]));
  AL_DFF_X al_97c00f94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[16]));
  AL_DFF_X al_e934978e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[17]));
  AL_DFF_X al_87fa5ea8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[18]));
  AL_DFF_X al_b2ae0585 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[1]));
  AL_DFF_X al_bd08f718 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[19]));
  AL_DFF_X al_285c24ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[20]));
  AL_DFF_X al_46fa2c51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[21]));
  AL_DFF_X al_dddffe66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[22]));
  AL_DFF_X al_69bcec30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[23]));
  AL_DFF_X al_763240af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[24]));
  AL_DFF_X al_382c5991 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[25]));
  AL_DFF_X al_ef23cd89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[26]));
  AL_DFF_X al_95153bad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[27]));
  AL_DFF_X al_e2f95295 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[28]));
  AL_DFF_X al_487aa1cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[2]));
  AL_DFF_X al_8f2192ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[29]));
  AL_DFF_X al_5d2c4aee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[30]));
  AL_DFF_X al_7dd1277d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[31]));
  AL_DFF_X al_865543c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[32]));
  AL_DFF_X al_76226423 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[33]));
  AL_DFF_X al_793fdde2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[34]));
  AL_DFF_X al_3cf133cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[35]));
  AL_DFF_X al_6a132b5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[36]));
  AL_DFF_X al_4bb00780 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[37]));
  AL_DFF_X al_60fe4490 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[38]));
  AL_DFF_X al_20c4a087 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[3]));
  AL_DFF_X al_5cba6296 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[39]));
  AL_DFF_X al_df767c75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[40]));
  AL_DFF_X al_90e55543 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[41]));
  AL_DFF_X al_d7831112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[42]));
  AL_DFF_X al_532d592f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[43]));
  AL_DFF_X al_4d99fc7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[44]));
  AL_DFF_X al_e21a95be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[45]));
  AL_DFF_X al_77bae67e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[46]));
  AL_DFF_X al_52aea47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e60d8647[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[47]));
  AL_DFF_X al_6f3b6f36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[4]));
  AL_DFF_X al_65441b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[5]));
  AL_DFF_X al_4520f572 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[6]));
  AL_DFF_X al_5c7979c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[7]));
  AL_DFF_X al_521f6b83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0f43754[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_86280a69[8]));
  AL_DFF_X al_8242878c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92faecea),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[0]));
  AL_DFF_X al_97cc8108 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[9]));
  AL_DFF_X al_dd844734 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[10]));
  AL_DFF_X al_2085b180 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[11]));
  AL_DFF_X al_af15f16b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[12]));
  AL_DFF_X al_b532d2b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[13]));
  AL_DFF_X al_24f342c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[14]));
  AL_DFF_X al_658b40a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[15]));
  AL_DFF_X al_1f0a38a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[16]));
  AL_DFF_X al_f73486ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[17]));
  AL_DFF_X al_d046aad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[18]));
  AL_DFF_X al_9db4ae72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[1]));
  AL_DFF_X al_b63781a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[19]));
  AL_DFF_X al_51a836e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[20]));
  AL_DFF_X al_548bc0a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[21]));
  AL_DFF_X al_7fa8fea5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[22]));
  AL_DFF_X al_52128586 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[23]));
  AL_DFF_X al_2db95c09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[2]));
  AL_DFF_X al_305166de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[3]));
  AL_DFF_X al_2b2258f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[4]));
  AL_DFF_X al_9ab8aa4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[5]));
  AL_DFF_X al_6e6df42a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[6]));
  AL_DFF_X al_3e314ca1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[7]));
  AL_DFF_X al_351935fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d3734717[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a4fb8f1[8]));
  AL_DFF_X al_d0db0ed5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e0dc7e9e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bade9fae[0]));
  AL_DFF_X al_b6b38c42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[22]));
  AL_DFF_X al_be28d7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[23]));
  AL_DFF_X al_32004ced (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[24]));
  AL_DFF_X al_6896cbd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[25]));
  AL_DFF_X al_dad9e5dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[26]));
  AL_DFF_X al_d95b8b3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[27]));
  AL_DFF_X al_48f1c0d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[28]));
  AL_DFF_X al_a7a7225e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[29]));
  AL_DFF_X al_e1bb2e8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[30]));
  AL_DFF_X al_e6ebb37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[31]));
  AL_DFF_X al_7ad3bce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[32]));
  AL_DFF_X al_61f89d90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[33]));
  AL_DFF_X al_89d161d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[34]));
  AL_DFF_X al_5bd6a5ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[35]));
  AL_DFF_X al_ca3356d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[36]));
  AL_DFF_X al_5180753c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[37]));
  AL_DFF_X al_eda4c4db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[38]));
  AL_DFF_X al_27995e9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[39]));
  AL_DFF_X al_29d6604e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[40]));
  AL_DFF_X al_fc116b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[41]));
  AL_DFF_X al_ecd40d74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[42]));
  AL_DFF_X al_e9f0bbd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[43]));
  AL_DFF_X al_1ce73241 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[44]));
  AL_DFF_X al_21d42456 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[45]));
  AL_DFF_X al_bdd6c687 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[46]));
  AL_DFF_X al_7f80953a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[47]));
  AL_DFF_X al_e27a616f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[48]));
  AL_DFF_X al_7ed39f7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[49]));
  AL_DFF_X al_a4351d0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[50]));
  AL_DFF_X al_6f8012d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[51]));
  AL_DFF_X al_5a326d2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[52]));
  AL_DFF_X al_93c5351f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3029c49a[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5181785e[53]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_111eec00 (
    .a(1'b0),
    .o({al_ddf49d7d,open_n86}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9f7e456f (
    .a(al_86280a69[23]),
    .b(al_3029c49a[23]),
    .c(al_ddf49d7d),
    .o({al_5613036,al_511419f7[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a3a84395 (
    .a(al_86280a69[24]),
    .b(al_3029c49a[24]),
    .c(al_5613036),
    .o({al_c86a97ab,al_511419f7[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7e919921 (
    .a(al_86280a69[25]),
    .b(al_3029c49a[25]),
    .c(al_c86a97ab),
    .o({al_ac57c034,al_511419f7[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_23f392e (
    .a(al_86280a69[26]),
    .b(al_3029c49a[26]),
    .c(al_ac57c034),
    .o({al_920c4e9a,al_511419f7[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6cde5deb (
    .a(al_86280a69[27]),
    .b(al_3029c49a[27]),
    .c(al_920c4e9a),
    .o({al_1283ff0b,al_511419f7[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_625156f9 (
    .a(al_86280a69[28]),
    .b(al_3029c49a[28]),
    .c(al_1283ff0b),
    .o({al_44359cb4,al_511419f7[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a01335c0 (
    .a(al_86280a69[29]),
    .b(al_3029c49a[29]),
    .c(al_44359cb4),
    .o({al_1fc8de48,al_511419f7[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f154b4a9 (
    .a(al_86280a69[30]),
    .b(al_3029c49a[30]),
    .c(al_1fc8de48),
    .o({al_9b620d8d,al_511419f7[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_992c8854 (
    .a(al_86280a69[31]),
    .b(al_3029c49a[31]),
    .c(al_9b620d8d),
    .o({al_c5542b59,al_511419f7[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_34d72715 (
    .a(al_86280a69[32]),
    .b(al_3029c49a[32]),
    .c(al_c5542b59),
    .o({al_fef84737,al_511419f7[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_be483d40 (
    .a(al_86280a69[33]),
    .b(al_3029c49a[33]),
    .c(al_fef84737),
    .o({al_d8cfcc23,al_511419f7[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b1e004c2 (
    .a(al_86280a69[34]),
    .b(al_3029c49a[34]),
    .c(al_d8cfcc23),
    .o({al_96385301,al_511419f7[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7af9ee70 (
    .a(al_86280a69[35]),
    .b(al_3029c49a[35]),
    .c(al_96385301),
    .o({al_2021f859,al_511419f7[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b8388692 (
    .a(al_86280a69[36]),
    .b(al_3029c49a[36]),
    .c(al_2021f859),
    .o({al_86a4ed5a,al_511419f7[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_66177baa (
    .a(al_86280a69[37]),
    .b(al_3029c49a[37]),
    .c(al_86a4ed5a),
    .o({al_52f700f5,al_511419f7[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f357a0b8 (
    .a(al_86280a69[38]),
    .b(al_3029c49a[38]),
    .c(al_52f700f5),
    .o({al_1024eced,al_511419f7[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_685f1a6a (
    .a(al_86280a69[39]),
    .b(al_3029c49a[39]),
    .c(al_1024eced),
    .o({al_55cc2fd4,al_511419f7[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1da79475 (
    .a(al_86280a69[40]),
    .b(al_3029c49a[40]),
    .c(al_55cc2fd4),
    .o({al_58146106,al_511419f7[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fe25ff10 (
    .a(al_86280a69[41]),
    .b(al_3029c49a[41]),
    .c(al_58146106),
    .o({al_b0f0b903,al_511419f7[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_96bdbfb4 (
    .a(al_86280a69[42]),
    .b(al_3029c49a[42]),
    .c(al_b0f0b903),
    .o({al_f01ea45c,al_511419f7[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d080bf03 (
    .a(al_86280a69[43]),
    .b(al_3029c49a[43]),
    .c(al_f01ea45c),
    .o({al_2b0b3830,al_511419f7[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc6624f3 (
    .a(al_86280a69[44]),
    .b(al_3029c49a[44]),
    .c(al_2b0b3830),
    .o({al_cc9bf94,al_511419f7[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8b85bedc (
    .a(al_86280a69[45]),
    .b(al_3029c49a[45]),
    .c(al_cc9bf94),
    .o({al_4a3ef4b7,al_511419f7[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_478886a0 (
    .a(al_86280a69[46]),
    .b(al_3029c49a[46]),
    .c(al_4a3ef4b7),
    .o({al_168ee139,al_511419f7[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_80d08431 (
    .a(al_86280a69[47]),
    .b(al_3029c49a[47]),
    .c(al_168ee139),
    .o({al_c52a2c84,al_511419f7[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_88f28a4c (
    .c(al_c52a2c84),
    .o({open_n89,al_511419f7[25]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_4cef2c6f (
    .a(al_3029c49a[50]),
    .b(al_3029c49a[51]),
    .c(al_3029c49a[52]),
    .d(al_3029c49a[53]),
    .e(al_3029c49a[54]),
    .f(al_511419f7[25]),
    .o(al_3a745b61));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    al_99a53fea (
    .a(al_3a745b61),
    .b(al_3029c49a[48]),
    .c(al_3029c49a[49]),
    .o(al_328e2c2d));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d6da71e (
    .a(al_328e2c2d),
    .b(al_86280a69[23]),
    .c(al_511419f7[0]),
    .o(al_f78b30ce[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1675244a (
    .a(al_328e2c2d),
    .b(al_86280a69[24]),
    .c(al_511419f7[1]),
    .o(al_f78b30ce[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_98f73b9d (
    .a(al_328e2c2d),
    .b(al_86280a69[25]),
    .c(al_511419f7[2]),
    .o(al_f78b30ce[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dca85609 (
    .a(al_328e2c2d),
    .b(al_86280a69[26]),
    .c(al_511419f7[3]),
    .o(al_f78b30ce[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d67ab856 (
    .a(al_328e2c2d),
    .b(al_86280a69[27]),
    .c(al_511419f7[4]),
    .o(al_f78b30ce[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_719b035e (
    .a(al_328e2c2d),
    .b(al_86280a69[28]),
    .c(al_511419f7[5]),
    .o(al_f78b30ce[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6e91bee6 (
    .a(al_328e2c2d),
    .b(al_86280a69[29]),
    .c(al_511419f7[6]),
    .o(al_f78b30ce[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d2e82af9 (
    .a(al_328e2c2d),
    .b(al_86280a69[30]),
    .c(al_511419f7[7]),
    .o(al_f78b30ce[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2e90ef1b (
    .a(al_328e2c2d),
    .b(al_86280a69[31]),
    .c(al_511419f7[8]),
    .o(al_f78b30ce[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1ba31507 (
    .a(al_328e2c2d),
    .b(al_86280a69[32]),
    .c(al_511419f7[9]),
    .o(al_f78b30ce[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e3a24f48 (
    .a(al_328e2c2d),
    .b(al_86280a69[33]),
    .c(al_511419f7[10]),
    .o(al_f78b30ce[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_877fa214 (
    .a(al_328e2c2d),
    .b(al_86280a69[34]),
    .c(al_511419f7[11]),
    .o(al_f78b30ce[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_94a24435 (
    .a(al_328e2c2d),
    .b(al_86280a69[35]),
    .c(al_511419f7[12]),
    .o(al_f78b30ce[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ad4e014b (
    .a(al_328e2c2d),
    .b(al_86280a69[36]),
    .c(al_511419f7[13]),
    .o(al_f78b30ce[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_28c6171d (
    .a(al_328e2c2d),
    .b(al_86280a69[37]),
    .c(al_511419f7[14]),
    .o(al_f78b30ce[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e9819304 (
    .a(al_328e2c2d),
    .b(al_86280a69[38]),
    .c(al_511419f7[15]),
    .o(al_f78b30ce[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5ffac473 (
    .a(al_328e2c2d),
    .b(al_86280a69[39]),
    .c(al_511419f7[16]),
    .o(al_f78b30ce[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f6cb0501 (
    .a(al_328e2c2d),
    .b(al_86280a69[40]),
    .c(al_511419f7[17]),
    .o(al_f78b30ce[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a125ed82 (
    .a(al_328e2c2d),
    .b(al_86280a69[41]),
    .c(al_511419f7[18]),
    .o(al_f78b30ce[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a0cbc027 (
    .a(al_328e2c2d),
    .b(al_86280a69[42]),
    .c(al_511419f7[19]),
    .o(al_f78b30ce[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8d129126 (
    .a(al_328e2c2d),
    .b(al_86280a69[43]),
    .c(al_511419f7[20]),
    .o(al_f78b30ce[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2ddffe9d (
    .a(al_328e2c2d),
    .b(al_86280a69[44]),
    .c(al_511419f7[21]),
    .o(al_f78b30ce[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e4011775 (
    .a(al_328e2c2d),
    .b(al_86280a69[45]),
    .c(al_511419f7[22]),
    .o(al_f78b30ce[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ef21c776 (
    .a(al_328e2c2d),
    .b(al_86280a69[46]),
    .c(al_511419f7[23]),
    .o(al_f78b30ce[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9d3d088e (
    .a(al_328e2c2d),
    .b(al_86280a69[47]),
    .c(al_511419f7[24]),
    .o(al_f78b30ce[47]));
  AL_DFF_X al_778492d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[0]));
  AL_DFF_X al_8f3b3f0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[9]));
  AL_DFF_X al_47b8f4e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[10]));
  AL_DFF_X al_8845c5ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[11]));
  AL_DFF_X al_5fc864fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[12]));
  AL_DFF_X al_a0dc2623 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[13]));
  AL_DFF_X al_761bd9d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[14]));
  AL_DFF_X al_b9327e5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[15]));
  AL_DFF_X al_676dcb26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[16]));
  AL_DFF_X al_ad454bcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[17]));
  AL_DFF_X al_f0cf5bc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[18]));
  AL_DFF_X al_78ac4ba6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[1]));
  AL_DFF_X al_3ffde316 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[19]));
  AL_DFF_X al_d092c16a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[20]));
  AL_DFF_X al_1001fa19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[21]));
  AL_DFF_X al_338154fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[22]));
  AL_DFF_X al_c88b5885 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[23]));
  AL_DFF_X al_30bd26c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[24]));
  AL_DFF_X al_b7b1c550 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[25]));
  AL_DFF_X al_1ca4837c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[26]));
  AL_DFF_X al_2e527677 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[27]));
  AL_DFF_X al_298b7369 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[28]));
  AL_DFF_X al_ca298abd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[2]));
  AL_DFF_X al_caf8e138 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[29]));
  AL_DFF_X al_ec9c69a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[30]));
  AL_DFF_X al_4361578e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[31]));
  AL_DFF_X al_fa96f76f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[32]));
  AL_DFF_X al_e6df4dda (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[33]));
  AL_DFF_X al_c64ee38d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[34]));
  AL_DFF_X al_a801e7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[35]));
  AL_DFF_X al_29aa3aef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[36]));
  AL_DFF_X al_71f8e79b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[37]));
  AL_DFF_X al_752d57b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[38]));
  AL_DFF_X al_e4d513eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[3]));
  AL_DFF_X al_f7c1bc89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[39]));
  AL_DFF_X al_c0e6fe3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[40]));
  AL_DFF_X al_f317df49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[41]));
  AL_DFF_X al_4695d973 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[42]));
  AL_DFF_X al_9a2fff89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[43]));
  AL_DFF_X al_1e1fc16d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[44]));
  AL_DFF_X al_23e7217 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[45]));
  AL_DFF_X al_3f3d6ed0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[46]));
  AL_DFF_X al_156ede5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f78b30ce[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[47]));
  AL_DFF_X al_31561449 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[4]));
  AL_DFF_X al_3a820202 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[5]));
  AL_DFF_X al_ffd2ced8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[6]));
  AL_DFF_X al_57781ea4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[7]));
  AL_DFF_X al_bf738445 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_86280a69[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9e3033a4[8]));
  AL_DFF_X al_10aaf554 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_328e2c2d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[0]));
  AL_DFF_X al_1d718554 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[9]));
  AL_DFF_X al_6a28bdfb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[10]));
  AL_DFF_X al_7cdf6eb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[11]));
  AL_DFF_X al_b76ae3f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[12]));
  AL_DFF_X al_386cef03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[13]));
  AL_DFF_X al_6828b3cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[14]));
  AL_DFF_X al_65943c5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[15]));
  AL_DFF_X al_6a3dba89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[16]));
  AL_DFF_X al_ea39b6a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[17]));
  AL_DFF_X al_6a04d929 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[18]));
  AL_DFF_X al_88e542eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[1]));
  AL_DFF_X al_6db50fc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[19]));
  AL_DFF_X al_1309af6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[20]));
  AL_DFF_X al_69ea4806 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[21]));
  AL_DFF_X al_a00d348a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[22]));
  AL_DFF_X al_e4df647b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[23]));
  AL_DFF_X al_e7071545 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[24]));
  AL_DFF_X al_80e576d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[2]));
  AL_DFF_X al_a573a023 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[3]));
  AL_DFF_X al_212b3e3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[4]));
  AL_DFF_X al_bd23b8c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[5]));
  AL_DFF_X al_bc676c36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[6]));
  AL_DFF_X al_2bfbe08e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[7]));
  AL_DFF_X al_a0bbcbb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a4fb8f1[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28f9bf01[8]));
  AL_DFF_X al_731835e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bade9fae[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f9ab06[0]));
  AL_DFF_X al_4c8b6992 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[21]));
  AL_DFF_X al_6894a2c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[22]));
  AL_DFF_X al_88037795 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[23]));
  AL_DFF_X al_1c043e35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[24]));
  AL_DFF_X al_8abd6ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[25]));
  AL_DFF_X al_8903232e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[26]));
  AL_DFF_X al_9bbc4f42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[27]));
  AL_DFF_X al_b5b64380 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[28]));
  AL_DFF_X al_5fb1c3cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[29]));
  AL_DFF_X al_765ac0c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[30]));
  AL_DFF_X al_2546c155 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[31]));
  AL_DFF_X al_58917b5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[32]));
  AL_DFF_X al_ed65ee59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[33]));
  AL_DFF_X al_fa25c375 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[34]));
  AL_DFF_X al_1788a3f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[35]));
  AL_DFF_X al_78c54952 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[36]));
  AL_DFF_X al_2a45d7fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[37]));
  AL_DFF_X al_11e68f2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[38]));
  AL_DFF_X al_f0b30116 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[39]));
  AL_DFF_X al_29bc3dbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[40]));
  AL_DFF_X al_45d785f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[41]));
  AL_DFF_X al_e7182a89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[42]));
  AL_DFF_X al_e18e3bd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[43]));
  AL_DFF_X al_373eea4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[44]));
  AL_DFF_X al_2584a47f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[45]));
  AL_DFF_X al_3ddcf3ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[46]));
  AL_DFF_X al_e4c202c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[47]));
  AL_DFF_X al_c82b8e48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[48]));
  AL_DFF_X al_3ae97dc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[49]));
  AL_DFF_X al_294e6dbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[50]));
  AL_DFF_X al_6a57a815 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[51]));
  AL_DFF_X al_9bf17f5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5181785e[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6a56028d[52]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_92d7cfc9 (
    .a(1'b0),
    .o({al_86e77cd0,open_n92}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_78c94b9f (
    .a(al_9e3033a4[22]),
    .b(al_5181785e[22]),
    .c(al_86e77cd0),
    .o({al_8b31527f,al_693e712c[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e407961a (
    .a(al_9e3033a4[23]),
    .b(al_5181785e[23]),
    .c(al_8b31527f),
    .o({al_1119be30,al_693e712c[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_15b3caf7 (
    .a(al_9e3033a4[24]),
    .b(al_5181785e[24]),
    .c(al_1119be30),
    .o({al_71939d74,al_693e712c[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2e3b1b6f (
    .a(al_9e3033a4[25]),
    .b(al_5181785e[25]),
    .c(al_71939d74),
    .o({al_d3344326,al_693e712c[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8a133eff (
    .a(al_9e3033a4[26]),
    .b(al_5181785e[26]),
    .c(al_d3344326),
    .o({al_e466bfff,al_693e712c[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9ef48331 (
    .a(al_9e3033a4[27]),
    .b(al_5181785e[27]),
    .c(al_e466bfff),
    .o({al_fe06d9ee,al_693e712c[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e7c6df3d (
    .a(al_9e3033a4[28]),
    .b(al_5181785e[28]),
    .c(al_fe06d9ee),
    .o({al_79cadb17,al_693e712c[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a7137e56 (
    .a(al_9e3033a4[29]),
    .b(al_5181785e[29]),
    .c(al_79cadb17),
    .o({al_e2799097,al_693e712c[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e700fbde (
    .a(al_9e3033a4[30]),
    .b(al_5181785e[30]),
    .c(al_e2799097),
    .o({al_12391d73,al_693e712c[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eaebd46e (
    .a(al_9e3033a4[31]),
    .b(al_5181785e[31]),
    .c(al_12391d73),
    .o({al_e4135f97,al_693e712c[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_46c530a6 (
    .a(al_9e3033a4[32]),
    .b(al_5181785e[32]),
    .c(al_e4135f97),
    .o({al_7c91f33c,al_693e712c[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d23a2e6 (
    .a(al_9e3033a4[33]),
    .b(al_5181785e[33]),
    .c(al_7c91f33c),
    .o({al_5576ac23,al_693e712c[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8ba0f402 (
    .a(al_9e3033a4[34]),
    .b(al_5181785e[34]),
    .c(al_5576ac23),
    .o({al_3f791172,al_693e712c[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2bf29f5d (
    .a(al_9e3033a4[35]),
    .b(al_5181785e[35]),
    .c(al_3f791172),
    .o({al_1c1093cd,al_693e712c[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_377f6a64 (
    .a(al_9e3033a4[36]),
    .b(al_5181785e[36]),
    .c(al_1c1093cd),
    .o({al_61436e1a,al_693e712c[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c2747c37 (
    .a(al_9e3033a4[37]),
    .b(al_5181785e[37]),
    .c(al_61436e1a),
    .o({al_bedba12b,al_693e712c[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a57f89a3 (
    .a(al_9e3033a4[38]),
    .b(al_5181785e[38]),
    .c(al_bedba12b),
    .o({al_c3463f35,al_693e712c[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_52503276 (
    .a(al_9e3033a4[39]),
    .b(al_5181785e[39]),
    .c(al_c3463f35),
    .o({al_fa3d49c2,al_693e712c[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_36210304 (
    .a(al_9e3033a4[40]),
    .b(al_5181785e[40]),
    .c(al_fa3d49c2),
    .o({al_caf86cb,al_693e712c[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_83b2c187 (
    .a(al_9e3033a4[41]),
    .b(al_5181785e[41]),
    .c(al_caf86cb),
    .o({al_603373a4,al_693e712c[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7f9cc07d (
    .a(al_9e3033a4[42]),
    .b(al_5181785e[42]),
    .c(al_603373a4),
    .o({al_236d63a,al_693e712c[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9815aad0 (
    .a(al_9e3033a4[43]),
    .b(al_5181785e[43]),
    .c(al_236d63a),
    .o({al_1e576ba8,al_693e712c[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d9f3f288 (
    .a(al_9e3033a4[44]),
    .b(al_5181785e[44]),
    .c(al_1e576ba8),
    .o({al_79f81494,al_693e712c[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c06bf399 (
    .a(al_9e3033a4[45]),
    .b(al_5181785e[45]),
    .c(al_79f81494),
    .o({al_921bd39c,al_693e712c[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6cca79cc (
    .a(al_9e3033a4[46]),
    .b(al_5181785e[46]),
    .c(al_921bd39c),
    .o({al_38de2714,al_693e712c[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ece11dcc (
    .a(al_9e3033a4[47]),
    .b(al_5181785e[47]),
    .c(al_38de2714),
    .o({al_b7b5bdbe,al_693e712c[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ac126b3a (
    .c(al_b7b5bdbe),
    .o({open_n95,al_693e712c[26]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fd13da36 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[22]),
    .c(al_693e712c[0]),
    .o(al_63579c4c[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d4e2464d (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[23]),
    .c(al_693e712c[1]),
    .o(al_63579c4c[23]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_dd9e78f6 (
    .a(al_5181785e[48]),
    .b(al_5181785e[49]),
    .c(al_5181785e[50]),
    .d(al_5181785e[51]),
    .e(al_5181785e[52]),
    .f(al_5181785e[53]),
    .o(al_43e60c58));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_9f8057ca (
    .a(al_43e60c58),
    .b(al_693e712c[26]),
    .o(al_d7aedbc5));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_69572de3 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[24]),
    .c(al_693e712c[2]),
    .o(al_63579c4c[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2e98e59f (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[25]),
    .c(al_693e712c[3]),
    .o(al_63579c4c[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ef05e4ac (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[26]),
    .c(al_693e712c[4]),
    .o(al_63579c4c[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7f79dde4 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[27]),
    .c(al_693e712c[5]),
    .o(al_63579c4c[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2b64b4b0 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[28]),
    .c(al_693e712c[6]),
    .o(al_63579c4c[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1a90d49b (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[29]),
    .c(al_693e712c[7]),
    .o(al_63579c4c[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6e9d85ca (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[30]),
    .c(al_693e712c[8]),
    .o(al_63579c4c[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bae6af86 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[31]),
    .c(al_693e712c[9]),
    .o(al_63579c4c[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5d402b23 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[32]),
    .c(al_693e712c[10]),
    .o(al_63579c4c[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3837e223 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[33]),
    .c(al_693e712c[11]),
    .o(al_63579c4c[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6d723816 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[34]),
    .c(al_693e712c[12]),
    .o(al_63579c4c[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cff8528f (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[35]),
    .c(al_693e712c[13]),
    .o(al_63579c4c[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8c07f325 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[36]),
    .c(al_693e712c[14]),
    .o(al_63579c4c[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ff60668 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[37]),
    .c(al_693e712c[15]),
    .o(al_63579c4c[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3541ed31 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[38]),
    .c(al_693e712c[16]),
    .o(al_63579c4c[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5be39203 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[39]),
    .c(al_693e712c[17]),
    .o(al_63579c4c[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_520a86fb (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[40]),
    .c(al_693e712c[18]),
    .o(al_63579c4c[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_29c43220 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[41]),
    .c(al_693e712c[19]),
    .o(al_63579c4c[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_66537c9b (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[42]),
    .c(al_693e712c[20]),
    .o(al_63579c4c[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_17cdb504 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[43]),
    .c(al_693e712c[21]),
    .o(al_63579c4c[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_233435dd (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[44]),
    .c(al_693e712c[22]),
    .o(al_63579c4c[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_93e12ef2 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[45]),
    .c(al_693e712c[23]),
    .o(al_63579c4c[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_66d747e (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[46]),
    .c(al_693e712c[24]),
    .o(al_63579c4c[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8500d919 (
    .a(al_d7aedbc5),
    .b(al_9e3033a4[47]),
    .c(al_693e712c[25]),
    .o(al_63579c4c[47]));
  AL_DFF_X al_f3cd9adc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[0]));
  AL_DFF_X al_e7ea96ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[9]));
  AL_DFF_X al_e60a4b75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[10]));
  AL_DFF_X al_768c89db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[11]));
  AL_DFF_X al_577d5734 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[12]));
  AL_DFF_X al_a99f0be7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[13]));
  AL_DFF_X al_4c433f58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[14]));
  AL_DFF_X al_2480314e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[15]));
  AL_DFF_X al_b356d127 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[16]));
  AL_DFF_X al_4bed32d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[17]));
  AL_DFF_X al_bf02b8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[18]));
  AL_DFF_X al_32a024f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[1]));
  AL_DFF_X al_63b7f535 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[19]));
  AL_DFF_X al_d8daba29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[20]));
  AL_DFF_X al_59297e7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[21]));
  AL_DFF_X al_a8879745 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[22]));
  AL_DFF_X al_2e37e242 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[23]));
  AL_DFF_X al_68ecfad4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[24]));
  AL_DFF_X al_c5c624a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[25]));
  AL_DFF_X al_6f972afa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[26]));
  AL_DFF_X al_bc6aa9c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[27]));
  AL_DFF_X al_5155a8cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[28]));
  AL_DFF_X al_15731b52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[2]));
  AL_DFF_X al_8344e864 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[29]));
  AL_DFF_X al_d8adada3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[30]));
  AL_DFF_X al_294d07bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[31]));
  AL_DFF_X al_d204c734 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[32]));
  AL_DFF_X al_9bb62962 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[33]));
  AL_DFF_X al_1a3044f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[34]));
  AL_DFF_X al_3bb92057 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[35]));
  AL_DFF_X al_2378c5e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[36]));
  AL_DFF_X al_85044b0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[37]));
  AL_DFF_X al_6e29154 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[38]));
  AL_DFF_X al_cef435d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[3]));
  AL_DFF_X al_ee1cc7b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[39]));
  AL_DFF_X al_be058005 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[40]));
  AL_DFF_X al_e775c22a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[41]));
  AL_DFF_X al_7fb473f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[42]));
  AL_DFF_X al_b18ce4b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[43]));
  AL_DFF_X al_4f51fe33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[44]));
  AL_DFF_X al_62b9ff43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[45]));
  AL_DFF_X al_e31a50ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[46]));
  AL_DFF_X al_cc010f62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_63579c4c[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[47]));
  AL_DFF_X al_cfd5f554 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[4]));
  AL_DFF_X al_1d00d0ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[5]));
  AL_DFF_X al_55f37d50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[6]));
  AL_DFF_X al_8c359765 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[7]));
  AL_DFF_X al_3ef03161 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e3033a4[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7397600a[8]));
  AL_DFF_X al_c3d38de3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d7aedbc5),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[0]));
  AL_DFF_X al_923b8b7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[9]));
  AL_DFF_X al_169f1f4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[10]));
  AL_DFF_X al_efa9cf81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[11]));
  AL_DFF_X al_40347cac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[12]));
  AL_DFF_X al_7e62cd04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[13]));
  AL_DFF_X al_522ff7f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[14]));
  AL_DFF_X al_1ec9927f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[15]));
  AL_DFF_X al_8da5b27f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[16]));
  AL_DFF_X al_1940b0c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[17]));
  AL_DFF_X al_9963f2cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[18]));
  AL_DFF_X al_8300be96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[1]));
  AL_DFF_X al_29de35dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[19]));
  AL_DFF_X al_72df9113 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[20]));
  AL_DFF_X al_9a9fe845 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[21]));
  AL_DFF_X al_3419f569 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[22]));
  AL_DFF_X al_bb18e908 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[23]));
  AL_DFF_X al_1ab353cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[24]));
  AL_DFF_X al_25e9d150 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[25]));
  AL_DFF_X al_fdde9169 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[2]));
  AL_DFF_X al_8ed6fff7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[3]));
  AL_DFF_X al_87ceead0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[4]));
  AL_DFF_X al_82ba71ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[5]));
  AL_DFF_X al_1d8cda8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[6]));
  AL_DFF_X al_f5a24378 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[7]));
  AL_DFF_X al_447b99fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28f9bf01[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c0ef3ebf[8]));
  AL_DFF_X al_c80db014 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8f9ab06[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fee4bd37[0]));
  AL_DFF_X al_633f3c75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[20]));
  AL_DFF_X al_30580cab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[21]));
  AL_DFF_X al_95d5352f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[22]));
  AL_DFF_X al_3b47431d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[23]));
  AL_DFF_X al_c7e09225 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[24]));
  AL_DFF_X al_a8119c77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[25]));
  AL_DFF_X al_b810a6a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[26]));
  AL_DFF_X al_158d721f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[27]));
  AL_DFF_X al_3e8afa31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[28]));
  AL_DFF_X al_318fb7a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[29]));
  AL_DFF_X al_787baa90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[30]));
  AL_DFF_X al_e2f518d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[31]));
  AL_DFF_X al_afc1eaf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[32]));
  AL_DFF_X al_e7830d04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[33]));
  AL_DFF_X al_c535209c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[34]));
  AL_DFF_X al_aaa7c793 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[35]));
  AL_DFF_X al_88990814 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[36]));
  AL_DFF_X al_9220a371 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[37]));
  AL_DFF_X al_992a20ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[38]));
  AL_DFF_X al_299638bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[39]));
  AL_DFF_X al_e7fea756 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[40]));
  AL_DFF_X al_42969552 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[41]));
  AL_DFF_X al_a0d101f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[42]));
  AL_DFF_X al_42aab558 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[43]));
  AL_DFF_X al_775df54f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[44]));
  AL_DFF_X al_5a04b285 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[45]));
  AL_DFF_X al_8fbfe2a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[46]));
  AL_DFF_X al_7f8d14bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[47]));
  AL_DFF_X al_416fd225 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[48]));
  AL_DFF_X al_aa83e995 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[49]));
  AL_DFF_X al_2263d8de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[50]));
  AL_DFF_X al_8010657e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a56028d[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6768e55[51]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_ddc7196a (
    .a(1'b0),
    .o({al_f67fc030,open_n98}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_decdcd1b (
    .a(al_7397600a[21]),
    .b(al_6a56028d[21]),
    .c(al_f67fc030),
    .o({al_e1b1f9c7,al_cabe3087[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_12a73ac1 (
    .a(al_7397600a[22]),
    .b(al_6a56028d[22]),
    .c(al_e1b1f9c7),
    .o({al_d27a6f7e,al_cabe3087[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ae7e7315 (
    .a(al_7397600a[23]),
    .b(al_6a56028d[23]),
    .c(al_d27a6f7e),
    .o({al_7932b374,al_cabe3087[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f6b2662c (
    .a(al_7397600a[24]),
    .b(al_6a56028d[24]),
    .c(al_7932b374),
    .o({al_93343d44,al_cabe3087[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_579211b2 (
    .a(al_7397600a[25]),
    .b(al_6a56028d[25]),
    .c(al_93343d44),
    .o({al_563f66f8,al_cabe3087[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_62138bf4 (
    .a(al_7397600a[26]),
    .b(al_6a56028d[26]),
    .c(al_563f66f8),
    .o({al_eb1ae9e7,al_cabe3087[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4a4fef62 (
    .a(al_7397600a[27]),
    .b(al_6a56028d[27]),
    .c(al_eb1ae9e7),
    .o({al_e483a091,al_cabe3087[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d679a9da (
    .a(al_7397600a[28]),
    .b(al_6a56028d[28]),
    .c(al_e483a091),
    .o({al_c3dfa0bb,al_cabe3087[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_781df829 (
    .a(al_7397600a[29]),
    .b(al_6a56028d[29]),
    .c(al_c3dfa0bb),
    .o({al_f67f9b7,al_cabe3087[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b4870139 (
    .a(al_7397600a[30]),
    .b(al_6a56028d[30]),
    .c(al_f67f9b7),
    .o({al_a6e65c64,al_cabe3087[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b61e70ff (
    .a(al_7397600a[31]),
    .b(al_6a56028d[31]),
    .c(al_a6e65c64),
    .o({al_a7b28424,al_cabe3087[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e2e18221 (
    .a(al_7397600a[32]),
    .b(al_6a56028d[32]),
    .c(al_a7b28424),
    .o({al_17c9f81e,al_cabe3087[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_378b7393 (
    .a(al_7397600a[33]),
    .b(al_6a56028d[33]),
    .c(al_17c9f81e),
    .o({al_ff089b0,al_cabe3087[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3fe638cf (
    .a(al_7397600a[34]),
    .b(al_6a56028d[34]),
    .c(al_ff089b0),
    .o({al_7f19c0cd,al_cabe3087[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e6bad64c (
    .a(al_7397600a[35]),
    .b(al_6a56028d[35]),
    .c(al_7f19c0cd),
    .o({al_aadee294,al_cabe3087[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_30f83fdb (
    .a(al_7397600a[36]),
    .b(al_6a56028d[36]),
    .c(al_aadee294),
    .o({al_1f32676d,al_cabe3087[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_41783706 (
    .a(al_7397600a[37]),
    .b(al_6a56028d[37]),
    .c(al_1f32676d),
    .o({al_e995362,al_cabe3087[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_966c63e4 (
    .a(al_7397600a[38]),
    .b(al_6a56028d[38]),
    .c(al_e995362),
    .o({al_28383266,al_cabe3087[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_12dd267a (
    .a(al_7397600a[39]),
    .b(al_6a56028d[39]),
    .c(al_28383266),
    .o({al_d33bf669,al_cabe3087[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_93f6b6f3 (
    .a(al_7397600a[40]),
    .b(al_6a56028d[40]),
    .c(al_d33bf669),
    .o({al_c70e8ffd,al_cabe3087[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2b0b5c9c (
    .a(al_7397600a[41]),
    .b(al_6a56028d[41]),
    .c(al_c70e8ffd),
    .o({al_f531391e,al_cabe3087[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_88c154c3 (
    .a(al_7397600a[42]),
    .b(al_6a56028d[42]),
    .c(al_f531391e),
    .o({al_c1cd2e91,al_cabe3087[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17de464e (
    .a(al_7397600a[43]),
    .b(al_6a56028d[43]),
    .c(al_c1cd2e91),
    .o({al_5361b136,al_cabe3087[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40de5145 (
    .a(al_7397600a[44]),
    .b(al_6a56028d[44]),
    .c(al_5361b136),
    .o({al_1f83c861,al_cabe3087[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_72d88331 (
    .a(al_7397600a[45]),
    .b(al_6a56028d[45]),
    .c(al_1f83c861),
    .o({al_1fd9ea3c,al_cabe3087[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_353be0aa (
    .a(al_7397600a[46]),
    .b(al_6a56028d[46]),
    .c(al_1fd9ea3c),
    .o({al_e10dc145,al_cabe3087[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c70ac8b2 (
    .a(al_7397600a[47]),
    .b(al_6a56028d[47]),
    .c(al_e10dc145),
    .o({al_dec1a002,al_cabe3087[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5a7aac85 (
    .c(al_dec1a002),
    .o({open_n101,al_cabe3087[27]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_285f8831 (
    .a(al_9e36993d),
    .b(al_7397600a[21]),
    .c(al_cabe3087[0]),
    .o(al_2c297489[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6034d936 (
    .a(al_9e36993d),
    .b(al_7397600a[22]),
    .c(al_cabe3087[1]),
    .o(al_2c297489[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f11b9504 (
    .a(al_9e36993d),
    .b(al_7397600a[23]),
    .c(al_cabe3087[2]),
    .o(al_2c297489[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e50e5e88 (
    .a(al_9e36993d),
    .b(al_7397600a[24]),
    .c(al_cabe3087[3]),
    .o(al_2c297489[24]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_948dbf8d (
    .a(al_6a56028d[48]),
    .b(al_6a56028d[49]),
    .c(al_6a56028d[50]),
    .d(al_6a56028d[51]),
    .e(al_6a56028d[52]),
    .f(al_cabe3087[27]),
    .o(al_9e36993d));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3c29dfb4 (
    .a(al_9e36993d),
    .b(al_7397600a[25]),
    .c(al_cabe3087[4]),
    .o(al_2c297489[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_be4fad80 (
    .a(al_9e36993d),
    .b(al_7397600a[26]),
    .c(al_cabe3087[5]),
    .o(al_2c297489[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d88731a4 (
    .a(al_9e36993d),
    .b(al_7397600a[27]),
    .c(al_cabe3087[6]),
    .o(al_2c297489[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2a8943 (
    .a(al_9e36993d),
    .b(al_7397600a[28]),
    .c(al_cabe3087[7]),
    .o(al_2c297489[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a1786b68 (
    .a(al_9e36993d),
    .b(al_7397600a[29]),
    .c(al_cabe3087[8]),
    .o(al_2c297489[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_93f2f040 (
    .a(al_9e36993d),
    .b(al_7397600a[30]),
    .c(al_cabe3087[9]),
    .o(al_2c297489[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_84afee8 (
    .a(al_9e36993d),
    .b(al_7397600a[31]),
    .c(al_cabe3087[10]),
    .o(al_2c297489[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_239e4fe5 (
    .a(al_9e36993d),
    .b(al_7397600a[32]),
    .c(al_cabe3087[11]),
    .o(al_2c297489[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fabbc6b0 (
    .a(al_9e36993d),
    .b(al_7397600a[33]),
    .c(al_cabe3087[12]),
    .o(al_2c297489[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_df5ed8a6 (
    .a(al_9e36993d),
    .b(al_7397600a[34]),
    .c(al_cabe3087[13]),
    .o(al_2c297489[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5cc71f85 (
    .a(al_9e36993d),
    .b(al_7397600a[35]),
    .c(al_cabe3087[14]),
    .o(al_2c297489[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_754717cb (
    .a(al_9e36993d),
    .b(al_7397600a[36]),
    .c(al_cabe3087[15]),
    .o(al_2c297489[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_329b827 (
    .a(al_9e36993d),
    .b(al_7397600a[37]),
    .c(al_cabe3087[16]),
    .o(al_2c297489[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_96ab2824 (
    .a(al_9e36993d),
    .b(al_7397600a[38]),
    .c(al_cabe3087[17]),
    .o(al_2c297489[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cbad0dd7 (
    .a(al_9e36993d),
    .b(al_7397600a[39]),
    .c(al_cabe3087[18]),
    .o(al_2c297489[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d9a0d7f6 (
    .a(al_9e36993d),
    .b(al_7397600a[40]),
    .c(al_cabe3087[19]),
    .o(al_2c297489[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c913391a (
    .a(al_9e36993d),
    .b(al_7397600a[41]),
    .c(al_cabe3087[20]),
    .o(al_2c297489[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_12ad321f (
    .a(al_9e36993d),
    .b(al_7397600a[42]),
    .c(al_cabe3087[21]),
    .o(al_2c297489[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_223e984 (
    .a(al_9e36993d),
    .b(al_7397600a[43]),
    .c(al_cabe3087[22]),
    .o(al_2c297489[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_89f1578d (
    .a(al_9e36993d),
    .b(al_7397600a[44]),
    .c(al_cabe3087[23]),
    .o(al_2c297489[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_45cf9b23 (
    .a(al_9e36993d),
    .b(al_7397600a[45]),
    .c(al_cabe3087[24]),
    .o(al_2c297489[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_beaeb7a (
    .a(al_9e36993d),
    .b(al_7397600a[46]),
    .c(al_cabe3087[25]),
    .o(al_2c297489[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_57be09b3 (
    .a(al_9e36993d),
    .b(al_7397600a[47]),
    .c(al_cabe3087[26]),
    .o(al_2c297489[47]));
  AL_DFF_X al_cda9996b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[0]));
  AL_DFF_X al_923ed742 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[9]));
  AL_DFF_X al_72a63ce9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[10]));
  AL_DFF_X al_80ca4007 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[11]));
  AL_DFF_X al_efdeba2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[12]));
  AL_DFF_X al_ec5df8e8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[13]));
  AL_DFF_X al_e817fdb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[14]));
  AL_DFF_X al_c240e7ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[15]));
  AL_DFF_X al_f1832113 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[16]));
  AL_DFF_X al_3bc1ae67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[17]));
  AL_DFF_X al_209800f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[18]));
  AL_DFF_X al_979a277f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[1]));
  AL_DFF_X al_46f2187d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[19]));
  AL_DFF_X al_b69cb58d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[20]));
  AL_DFF_X al_7aa0433e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[21]));
  AL_DFF_X al_403de344 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[22]));
  AL_DFF_X al_92964f61 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[23]));
  AL_DFF_X al_2671ab98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[24]));
  AL_DFF_X al_f7ea9ab4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[25]));
  AL_DFF_X al_f80a4e54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[26]));
  AL_DFF_X al_63820373 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[27]));
  AL_DFF_X al_cbfcf96d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[28]));
  AL_DFF_X al_765c24f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[2]));
  AL_DFF_X al_a244ec59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[29]));
  AL_DFF_X al_44e3cb3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[30]));
  AL_DFF_X al_2675f0c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[31]));
  AL_DFF_X al_84243159 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[32]));
  AL_DFF_X al_a6d496a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[33]));
  AL_DFF_X al_56d32acc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[34]));
  AL_DFF_X al_f236b1d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[35]));
  AL_DFF_X al_f5870913 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[36]));
  AL_DFF_X al_38412d5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[37]));
  AL_DFF_X al_76a9ab54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[38]));
  AL_DFF_X al_fb29211d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[3]));
  AL_DFF_X al_64c8f2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[39]));
  AL_DFF_X al_140f9ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[40]));
  AL_DFF_X al_804a7936 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[41]));
  AL_DFF_X al_495afcaa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[42]));
  AL_DFF_X al_aaec55f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[43]));
  AL_DFF_X al_ace07f3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[44]));
  AL_DFF_X al_1f30d006 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[45]));
  AL_DFF_X al_cbadc65b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[46]));
  AL_DFF_X al_3e64dc1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c297489[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[47]));
  AL_DFF_X al_491f86bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[4]));
  AL_DFF_X al_6581ed8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[5]));
  AL_DFF_X al_9181e10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[6]));
  AL_DFF_X al_8c9b73c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[7]));
  AL_DFF_X al_b09383db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7397600a[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e4be4089[8]));
  AL_DFF_X al_bd0add42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9e36993d),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[0]));
  AL_DFF_X al_ff093264 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[9]));
  AL_DFF_X al_eb6bd45d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[10]));
  AL_DFF_X al_205f9953 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[11]));
  AL_DFF_X al_960f7191 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[12]));
  AL_DFF_X al_f6d4da02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[13]));
  AL_DFF_X al_59bee5b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[14]));
  AL_DFF_X al_a8d52617 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[15]));
  AL_DFF_X al_18a61cf7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[16]));
  AL_DFF_X al_78c13320 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[17]));
  AL_DFF_X al_a3588029 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[18]));
  AL_DFF_X al_c14b0412 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[1]));
  AL_DFF_X al_f930372a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[19]));
  AL_DFF_X al_e6fc5803 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[20]));
  AL_DFF_X al_14e72213 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[21]));
  AL_DFF_X al_dfd0c72b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[22]));
  AL_DFF_X al_57aeb8b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[23]));
  AL_DFF_X al_dc949970 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[24]));
  AL_DFF_X al_55dcdd73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[25]));
  AL_DFF_X al_42d00463 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[26]));
  AL_DFF_X al_c7de715a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[2]));
  AL_DFF_X al_9b66f075 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[3]));
  AL_DFF_X al_28b9079f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[4]));
  AL_DFF_X al_35d72850 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[5]));
  AL_DFF_X al_1eeae453 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[6]));
  AL_DFF_X al_3df9f52e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[7]));
  AL_DFF_X al_d1a9be38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c0ef3ebf[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d71a2aba[8]));
  AL_DFF_X al_9f3702f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_fee4bd37[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e0e2aae4[0]));
  AL_DFF_X al_69b28580 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[19]));
  AL_DFF_X al_db91fd4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[20]));
  AL_DFF_X al_3ca62244 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[21]));
  AL_DFF_X al_5e7b6c06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[22]));
  AL_DFF_X al_e6e03be4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[23]));
  AL_DFF_X al_864ff74e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[24]));
  AL_DFF_X al_e32337ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[25]));
  AL_DFF_X al_415c82ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[26]));
  AL_DFF_X al_8f09bd6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[27]));
  AL_DFF_X al_82d25619 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[28]));
  AL_DFF_X al_b259398b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[29]));
  AL_DFF_X al_7c02a6e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[30]));
  AL_DFF_X al_8fef6922 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[31]));
  AL_DFF_X al_7605098b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[32]));
  AL_DFF_X al_fea73481 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[33]));
  AL_DFF_X al_3c5479a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[34]));
  AL_DFF_X al_4744276a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[35]));
  AL_DFF_X al_d2d734ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[36]));
  AL_DFF_X al_317af8a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[37]));
  AL_DFF_X al_ce4f0760 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[38]));
  AL_DFF_X al_a264ffec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[39]));
  AL_DFF_X al_eb7ce11c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[40]));
  AL_DFF_X al_9ba781a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[41]));
  AL_DFF_X al_a9ba82d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[42]));
  AL_DFF_X al_b2b01028 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[43]));
  AL_DFF_X al_eacb78ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[44]));
  AL_DFF_X al_fb4009b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[45]));
  AL_DFF_X al_d764358 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[46]));
  AL_DFF_X al_69b504ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[47]));
  AL_DFF_X al_85d87fee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[48]));
  AL_DFF_X al_d7833dc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[49]));
  AL_DFF_X al_c60b88d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6768e55[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_222a5f4d[50]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_1066ffed (
    .a(1'b0),
    .o({al_8302a2a2,open_n104}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d18b138b (
    .a(al_e4be4089[20]),
    .b(al_b6768e55[20]),
    .c(al_8302a2a2),
    .o({al_78579729,al_c307e46[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_86d29383 (
    .a(al_e4be4089[21]),
    .b(al_b6768e55[21]),
    .c(al_78579729),
    .o({al_cce3e61c,al_c307e46[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4fbe4ec1 (
    .a(al_e4be4089[22]),
    .b(al_b6768e55[22]),
    .c(al_cce3e61c),
    .o({al_edfe5545,al_c307e46[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2f64522e (
    .a(al_e4be4089[23]),
    .b(al_b6768e55[23]),
    .c(al_edfe5545),
    .o({al_8afadf84,al_c307e46[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cb781d3f (
    .a(al_e4be4089[24]),
    .b(al_b6768e55[24]),
    .c(al_8afadf84),
    .o({al_91c4f866,al_c307e46[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9fc0556f (
    .a(al_e4be4089[25]),
    .b(al_b6768e55[25]),
    .c(al_91c4f866),
    .o({al_dfb38e7,al_c307e46[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_afb51a7d (
    .a(al_e4be4089[26]),
    .b(al_b6768e55[26]),
    .c(al_dfb38e7),
    .o({al_ea5a8045,al_c307e46[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f1ac0c32 (
    .a(al_e4be4089[27]),
    .b(al_b6768e55[27]),
    .c(al_ea5a8045),
    .o({al_5594316d,al_c307e46[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dc85e8ae (
    .a(al_e4be4089[28]),
    .b(al_b6768e55[28]),
    .c(al_5594316d),
    .o({al_802edd1b,al_c307e46[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ac598961 (
    .a(al_e4be4089[29]),
    .b(al_b6768e55[29]),
    .c(al_802edd1b),
    .o({al_4ed141e3,al_c307e46[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ed754f07 (
    .a(al_e4be4089[30]),
    .b(al_b6768e55[30]),
    .c(al_4ed141e3),
    .o({al_a9bde1cf,al_c307e46[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_963dfd4e (
    .a(al_e4be4089[31]),
    .b(al_b6768e55[31]),
    .c(al_a9bde1cf),
    .o({al_b879dc6c,al_c307e46[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b4ac4718 (
    .a(al_e4be4089[32]),
    .b(al_b6768e55[32]),
    .c(al_b879dc6c),
    .o({al_8f601d11,al_c307e46[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1e378a63 (
    .a(al_e4be4089[33]),
    .b(al_b6768e55[33]),
    .c(al_8f601d11),
    .o({al_1861ccb9,al_c307e46[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_afd646a7 (
    .a(al_e4be4089[34]),
    .b(al_b6768e55[34]),
    .c(al_1861ccb9),
    .o({al_417b1b7f,al_c307e46[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d6ff6348 (
    .a(al_e4be4089[35]),
    .b(al_b6768e55[35]),
    .c(al_417b1b7f),
    .o({al_a4400d46,al_c307e46[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b743ef35 (
    .a(al_e4be4089[36]),
    .b(al_b6768e55[36]),
    .c(al_a4400d46),
    .o({al_59eab12e,al_c307e46[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_781e500f (
    .a(al_e4be4089[37]),
    .b(al_b6768e55[37]),
    .c(al_59eab12e),
    .o({al_1af64e4d,al_c307e46[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c2458f1c (
    .a(al_e4be4089[38]),
    .b(al_b6768e55[38]),
    .c(al_1af64e4d),
    .o({al_ecd39a7,al_c307e46[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f8c6621d (
    .a(al_e4be4089[39]),
    .b(al_b6768e55[39]),
    .c(al_ecd39a7),
    .o({al_a7d6fdcd,al_c307e46[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ebdbe3ff (
    .a(al_e4be4089[40]),
    .b(al_b6768e55[40]),
    .c(al_a7d6fdcd),
    .o({al_7de07321,al_c307e46[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc71dc1f (
    .a(al_e4be4089[41]),
    .b(al_b6768e55[41]),
    .c(al_7de07321),
    .o({al_df148873,al_c307e46[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f8e47c45 (
    .a(al_e4be4089[42]),
    .b(al_b6768e55[42]),
    .c(al_df148873),
    .o({al_1f49b9e4,al_c307e46[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cdafa0f3 (
    .a(al_e4be4089[43]),
    .b(al_b6768e55[43]),
    .c(al_1f49b9e4),
    .o({al_832fb3e,al_c307e46[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a0f4601c (
    .a(al_e4be4089[44]),
    .b(al_b6768e55[44]),
    .c(al_832fb3e),
    .o({al_2d137dff,al_c307e46[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_58d58286 (
    .a(al_e4be4089[45]),
    .b(al_b6768e55[45]),
    .c(al_2d137dff),
    .o({al_fd484a6d,al_c307e46[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_85bd46c1 (
    .a(al_e4be4089[46]),
    .b(al_b6768e55[46]),
    .c(al_fd484a6d),
    .o({al_1d7722f2,al_c307e46[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cb371cb (
    .a(al_e4be4089[47]),
    .b(al_b6768e55[47]),
    .c(al_1d7722f2),
    .o({al_83dc3e4f,al_c307e46[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4cdcc470 (
    .c(al_83dc3e4f),
    .o({open_n107,al_c307e46[28]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_812d1ca8 (
    .a(al_e7c4a377),
    .b(al_e4be4089[20]),
    .c(al_c307e46[0]),
    .o(al_9857f6b5[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ce868b8d (
    .a(al_e7c4a377),
    .b(al_e4be4089[21]),
    .c(al_c307e46[1]),
    .o(al_9857f6b5[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_34b7cb0f (
    .a(al_e7c4a377),
    .b(al_e4be4089[22]),
    .c(al_c307e46[2]),
    .o(al_9857f6b5[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_aeb1fe37 (
    .a(al_e7c4a377),
    .b(al_e4be4089[23]),
    .c(al_c307e46[3]),
    .o(al_9857f6b5[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_162fda05 (
    .a(al_e7c4a377),
    .b(al_e4be4089[24]),
    .c(al_c307e46[4]),
    .o(al_9857f6b5[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f0639d5d (
    .a(al_e7c4a377),
    .b(al_e4be4089[25]),
    .c(al_c307e46[5]),
    .o(al_9857f6b5[25]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_255f48b6 (
    .a(al_b6768e55[48]),
    .b(al_b6768e55[49]),
    .c(al_b6768e55[50]),
    .d(al_b6768e55[51]),
    .e(al_c307e46[28]),
    .o(al_e7c4a377));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ce09416f (
    .a(al_e7c4a377),
    .b(al_e4be4089[26]),
    .c(al_c307e46[6]),
    .o(al_9857f6b5[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dd419afc (
    .a(al_e7c4a377),
    .b(al_e4be4089[27]),
    .c(al_c307e46[7]),
    .o(al_9857f6b5[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2f3c91a (
    .a(al_e7c4a377),
    .b(al_e4be4089[28]),
    .c(al_c307e46[8]),
    .o(al_9857f6b5[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_601e8e7a (
    .a(al_e7c4a377),
    .b(al_e4be4089[29]),
    .c(al_c307e46[9]),
    .o(al_9857f6b5[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7ac0d4fa (
    .a(al_e7c4a377),
    .b(al_e4be4089[30]),
    .c(al_c307e46[10]),
    .o(al_9857f6b5[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_65aa7b93 (
    .a(al_e7c4a377),
    .b(al_e4be4089[31]),
    .c(al_c307e46[11]),
    .o(al_9857f6b5[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f0e1657c (
    .a(al_e7c4a377),
    .b(al_e4be4089[32]),
    .c(al_c307e46[12]),
    .o(al_9857f6b5[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c5435094 (
    .a(al_e7c4a377),
    .b(al_e4be4089[33]),
    .c(al_c307e46[13]),
    .o(al_9857f6b5[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_483f37ec (
    .a(al_e7c4a377),
    .b(al_e4be4089[34]),
    .c(al_c307e46[14]),
    .o(al_9857f6b5[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_16f38105 (
    .a(al_e7c4a377),
    .b(al_e4be4089[35]),
    .c(al_c307e46[15]),
    .o(al_9857f6b5[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b6e864b (
    .a(al_e7c4a377),
    .b(al_e4be4089[36]),
    .c(al_c307e46[16]),
    .o(al_9857f6b5[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a3be4e67 (
    .a(al_e7c4a377),
    .b(al_e4be4089[37]),
    .c(al_c307e46[17]),
    .o(al_9857f6b5[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_85a5011e (
    .a(al_e7c4a377),
    .b(al_e4be4089[38]),
    .c(al_c307e46[18]),
    .o(al_9857f6b5[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_88027cf6 (
    .a(al_e7c4a377),
    .b(al_e4be4089[39]),
    .c(al_c307e46[19]),
    .o(al_9857f6b5[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4f5ab8ed (
    .a(al_e7c4a377),
    .b(al_e4be4089[40]),
    .c(al_c307e46[20]),
    .o(al_9857f6b5[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7664ad16 (
    .a(al_e7c4a377),
    .b(al_e4be4089[41]),
    .c(al_c307e46[21]),
    .o(al_9857f6b5[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2da9d129 (
    .a(al_e7c4a377),
    .b(al_e4be4089[42]),
    .c(al_c307e46[22]),
    .o(al_9857f6b5[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2fd7b7ba (
    .a(al_e7c4a377),
    .b(al_e4be4089[43]),
    .c(al_c307e46[23]),
    .o(al_9857f6b5[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c5029e31 (
    .a(al_e7c4a377),
    .b(al_e4be4089[44]),
    .c(al_c307e46[24]),
    .o(al_9857f6b5[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_60f49d67 (
    .a(al_e7c4a377),
    .b(al_e4be4089[45]),
    .c(al_c307e46[25]),
    .o(al_9857f6b5[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d8370b5a (
    .a(al_e7c4a377),
    .b(al_e4be4089[46]),
    .c(al_c307e46[26]),
    .o(al_9857f6b5[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a84958cf (
    .a(al_e7c4a377),
    .b(al_e4be4089[47]),
    .c(al_c307e46[27]),
    .o(al_9857f6b5[47]));
  AL_DFF_X al_bf989e85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[0]));
  AL_DFF_X al_c8935819 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[9]));
  AL_DFF_X al_ebcdc75e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[10]));
  AL_DFF_X al_545e21b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[11]));
  AL_DFF_X al_bb96ab66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[12]));
  AL_DFF_X al_f118d545 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[13]));
  AL_DFF_X al_57da5d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[14]));
  AL_DFF_X al_f560c43d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[15]));
  AL_DFF_X al_aa97977e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[16]));
  AL_DFF_X al_fe7a2e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[17]));
  AL_DFF_X al_b9cc4686 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[18]));
  AL_DFF_X al_2e984074 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[1]));
  AL_DFF_X al_284c553d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[19]));
  AL_DFF_X al_ca9d183d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[20]));
  AL_DFF_X al_f0c80a71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[21]));
  AL_DFF_X al_ea209e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[22]));
  AL_DFF_X al_70fe1a65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[23]));
  AL_DFF_X al_2295ce21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[24]));
  AL_DFF_X al_1f1374ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[25]));
  AL_DFF_X al_6f3390bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[26]));
  AL_DFF_X al_f7a223fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[27]));
  AL_DFF_X al_c09df45f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[28]));
  AL_DFF_X al_535a9912 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[2]));
  AL_DFF_X al_3a93cf1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[29]));
  AL_DFF_X al_8faf18cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[30]));
  AL_DFF_X al_8d1169b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[31]));
  AL_DFF_X al_e598d9b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[32]));
  AL_DFF_X al_5b6c618f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[33]));
  AL_DFF_X al_f23c4574 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[34]));
  AL_DFF_X al_a2efe2a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[35]));
  AL_DFF_X al_b662ac3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[36]));
  AL_DFF_X al_41eb41f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[37]));
  AL_DFF_X al_46b2411e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[38]));
  AL_DFF_X al_f6ea2f86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[3]));
  AL_DFF_X al_e4f716e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[39]));
  AL_DFF_X al_f359d1b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[40]));
  AL_DFF_X al_30b32744 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[41]));
  AL_DFF_X al_a35fd891 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[42]));
  AL_DFF_X al_4f161ddc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[43]));
  AL_DFF_X al_febad3d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[44]));
  AL_DFF_X al_b52214c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[45]));
  AL_DFF_X al_607e7f0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[46]));
  AL_DFF_X al_bceeb4f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9857f6b5[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[47]));
  AL_DFF_X al_2e40cbdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[4]));
  AL_DFF_X al_e28d3f94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[5]));
  AL_DFF_X al_166eb818 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[6]));
  AL_DFF_X al_9ac0216c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[7]));
  AL_DFF_X al_34550309 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e4be4089[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4a463b38[8]));
  AL_DFF_X al_3225089f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7c4a377),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[0]));
  AL_DFF_X al_7819b3b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[9]));
  AL_DFF_X al_1dda5439 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[10]));
  AL_DFF_X al_3882f4c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[11]));
  AL_DFF_X al_655b5d8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[12]));
  AL_DFF_X al_f4b7f123 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[13]));
  AL_DFF_X al_47f6d32a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[14]));
  AL_DFF_X al_e1a12649 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[15]));
  AL_DFF_X al_3f8196dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[16]));
  AL_DFF_X al_ce2f65bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[17]));
  AL_DFF_X al_fa79b29c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[18]));
  AL_DFF_X al_73378a69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[1]));
  AL_DFF_X al_22207116 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[19]));
  AL_DFF_X al_bbcf803d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[20]));
  AL_DFF_X al_691d7225 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[21]));
  AL_DFF_X al_1c79d934 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[22]));
  AL_DFF_X al_2c5f7702 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[23]));
  AL_DFF_X al_6b2700b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[24]));
  AL_DFF_X al_33a442cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[25]));
  AL_DFF_X al_36b7a216 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[26]));
  AL_DFF_X al_24fe5cb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[27]));
  AL_DFF_X al_76e094a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[2]));
  AL_DFF_X al_a48fc827 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[3]));
  AL_DFF_X al_819f1f51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[4]));
  AL_DFF_X al_c0b8a80c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[5]));
  AL_DFF_X al_ab9d283e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[6]));
  AL_DFF_X al_75e5e297 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[7]));
  AL_DFF_X al_9220c6ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d71a2aba[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7a3cd65[8]));
  AL_DFF_X al_8f584f17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e0e2aae4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5db428bb[0]));
  AL_DFF_X al_ee2cb809 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[18]));
  AL_DFF_X al_34f73d8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[19]));
  AL_DFF_X al_62b83983 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[20]));
  AL_DFF_X al_331dd442 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[21]));
  AL_DFF_X al_e2af1298 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[22]));
  AL_DFF_X al_8cefc710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[23]));
  AL_DFF_X al_9e78ebe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[24]));
  AL_DFF_X al_e4dba65e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[25]));
  AL_DFF_X al_58dd9cd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[26]));
  AL_DFF_X al_58f5fe4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[27]));
  AL_DFF_X al_312c80d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[28]));
  AL_DFF_X al_e2488f31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[29]));
  AL_DFF_X al_4da471a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[30]));
  AL_DFF_X al_b8a48d7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[31]));
  AL_DFF_X al_abd1ce39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[32]));
  AL_DFF_X al_967e6603 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[33]));
  AL_DFF_X al_174d298e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[34]));
  AL_DFF_X al_8e25d438 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[35]));
  AL_DFF_X al_6099cc37 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[36]));
  AL_DFF_X al_c09f9a1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[37]));
  AL_DFF_X al_88981dfb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[38]));
  AL_DFF_X al_6e49947 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[39]));
  AL_DFF_X al_d4d5cde (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[40]));
  AL_DFF_X al_b6914311 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[41]));
  AL_DFF_X al_fa52c63b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[42]));
  AL_DFF_X al_2c912071 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[43]));
  AL_DFF_X al_485b6e90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[44]));
  AL_DFF_X al_c9eaba60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[45]));
  AL_DFF_X al_b8807642 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[46]));
  AL_DFF_X al_76ecf667 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[47]));
  AL_DFF_X al_5fed62a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[48]));
  AL_DFF_X al_484aa8f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_222a5f4d[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d1a07609[49]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_bd29075c (
    .a(1'b0),
    .o({al_153001b0,open_n110}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d19768f8 (
    .a(al_4a463b38[19]),
    .b(al_222a5f4d[19]),
    .c(al_153001b0),
    .o({al_90b73cc5,al_794ac8f[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4ab1d7f3 (
    .a(al_4a463b38[20]),
    .b(al_222a5f4d[20]),
    .c(al_90b73cc5),
    .o({al_6cc49207,al_794ac8f[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c7a400e3 (
    .a(al_4a463b38[21]),
    .b(al_222a5f4d[21]),
    .c(al_6cc49207),
    .o({al_88ebd806,al_794ac8f[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc06dcbd (
    .a(al_4a463b38[22]),
    .b(al_222a5f4d[22]),
    .c(al_88ebd806),
    .o({al_9ba3e8a0,al_794ac8f[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3b4b8008 (
    .a(al_4a463b38[23]),
    .b(al_222a5f4d[23]),
    .c(al_9ba3e8a0),
    .o({al_c1436409,al_794ac8f[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f6c08999 (
    .a(al_4a463b38[24]),
    .b(al_222a5f4d[24]),
    .c(al_c1436409),
    .o({al_a907358b,al_794ac8f[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_57901726 (
    .a(al_4a463b38[25]),
    .b(al_222a5f4d[25]),
    .c(al_a907358b),
    .o({al_7c92a6e7,al_794ac8f[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f20a6669 (
    .a(al_4a463b38[26]),
    .b(al_222a5f4d[26]),
    .c(al_7c92a6e7),
    .o({al_2848275b,al_794ac8f[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bf98e697 (
    .a(al_4a463b38[27]),
    .b(al_222a5f4d[27]),
    .c(al_2848275b),
    .o({al_1cb31d61,al_794ac8f[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a9605403 (
    .a(al_4a463b38[28]),
    .b(al_222a5f4d[28]),
    .c(al_1cb31d61),
    .o({al_ddf9bf5e,al_794ac8f[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eb68ded2 (
    .a(al_4a463b38[29]),
    .b(al_222a5f4d[29]),
    .c(al_ddf9bf5e),
    .o({al_4cef4276,al_794ac8f[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9d1fb8b8 (
    .a(al_4a463b38[30]),
    .b(al_222a5f4d[30]),
    .c(al_4cef4276),
    .o({al_6cf3b362,al_794ac8f[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dfb02c5a (
    .a(al_4a463b38[31]),
    .b(al_222a5f4d[31]),
    .c(al_6cf3b362),
    .o({al_e0b0ba1d,al_794ac8f[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_452ec2ef (
    .a(al_4a463b38[32]),
    .b(al_222a5f4d[32]),
    .c(al_e0b0ba1d),
    .o({al_5c52a055,al_794ac8f[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_72bf4675 (
    .a(al_4a463b38[33]),
    .b(al_222a5f4d[33]),
    .c(al_5c52a055),
    .o({al_90d0cde9,al_794ac8f[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_50653447 (
    .a(al_4a463b38[34]),
    .b(al_222a5f4d[34]),
    .c(al_90d0cde9),
    .o({al_b506c4,al_794ac8f[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b8f26dd (
    .a(al_4a463b38[35]),
    .b(al_222a5f4d[35]),
    .c(al_b506c4),
    .o({al_63ccb9ff,al_794ac8f[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_72f09045 (
    .a(al_4a463b38[36]),
    .b(al_222a5f4d[36]),
    .c(al_63ccb9ff),
    .o({al_72ec7913,al_794ac8f[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ef0ae947 (
    .a(al_4a463b38[37]),
    .b(al_222a5f4d[37]),
    .c(al_72ec7913),
    .o({al_a727e78e,al_794ac8f[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9d3bc524 (
    .a(al_4a463b38[38]),
    .b(al_222a5f4d[38]),
    .c(al_a727e78e),
    .o({al_61742d3d,al_794ac8f[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_aaeec10a (
    .a(al_4a463b38[39]),
    .b(al_222a5f4d[39]),
    .c(al_61742d3d),
    .o({al_da23077d,al_794ac8f[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a3e5c310 (
    .a(al_4a463b38[40]),
    .b(al_222a5f4d[40]),
    .c(al_da23077d),
    .o({al_d907d72,al_794ac8f[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f620c21 (
    .a(al_4a463b38[41]),
    .b(al_222a5f4d[41]),
    .c(al_d907d72),
    .o({al_941ec574,al_794ac8f[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6cb797d5 (
    .a(al_4a463b38[42]),
    .b(al_222a5f4d[42]),
    .c(al_941ec574),
    .o({al_e915b010,al_794ac8f[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_75d99e98 (
    .a(al_4a463b38[43]),
    .b(al_222a5f4d[43]),
    .c(al_e915b010),
    .o({al_4f44504e,al_794ac8f[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3728e305 (
    .a(al_4a463b38[44]),
    .b(al_222a5f4d[44]),
    .c(al_4f44504e),
    .o({al_30d605ba,al_794ac8f[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_db3a6775 (
    .a(al_4a463b38[45]),
    .b(al_222a5f4d[45]),
    .c(al_30d605ba),
    .o({al_8c151872,al_794ac8f[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_42ffdc1b (
    .a(al_4a463b38[46]),
    .b(al_222a5f4d[46]),
    .c(al_8c151872),
    .o({al_e2a656fd,al_794ac8f[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dce5e411 (
    .a(al_4a463b38[47]),
    .b(al_222a5f4d[47]),
    .c(al_e2a656fd),
    .o({al_55ab11c1,al_794ac8f[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_863c18e (
    .c(al_55ab11c1),
    .o({open_n113,al_794ac8f[29]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a97a84a2 (
    .a(al_281a7b5c),
    .b(al_4a463b38[19]),
    .c(al_794ac8f[0]),
    .o(al_e343d659[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9bc6d77a (
    .a(al_281a7b5c),
    .b(al_4a463b38[20]),
    .c(al_794ac8f[1]),
    .o(al_e343d659[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4fa5015c (
    .a(al_281a7b5c),
    .b(al_4a463b38[21]),
    .c(al_794ac8f[2]),
    .o(al_e343d659[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9447a0dd (
    .a(al_281a7b5c),
    .b(al_4a463b38[22]),
    .c(al_794ac8f[3]),
    .o(al_e343d659[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2cc9bd8 (
    .a(al_281a7b5c),
    .b(al_4a463b38[23]),
    .c(al_794ac8f[4]),
    .o(al_e343d659[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3b7b6b52 (
    .a(al_281a7b5c),
    .b(al_4a463b38[24]),
    .c(al_794ac8f[5]),
    .o(al_e343d659[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_67fe5ba4 (
    .a(al_281a7b5c),
    .b(al_4a463b38[25]),
    .c(al_794ac8f[6]),
    .o(al_e343d659[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1fa28c08 (
    .a(al_281a7b5c),
    .b(al_4a463b38[26]),
    .c(al_794ac8f[7]),
    .o(al_e343d659[26]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    al_8da17227 (
    .a(al_222a5f4d[48]),
    .b(al_222a5f4d[49]),
    .c(al_222a5f4d[50]),
    .d(al_794ac8f[29]),
    .o(al_281a7b5c));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fea31acc (
    .a(al_281a7b5c),
    .b(al_4a463b38[27]),
    .c(al_794ac8f[8]),
    .o(al_e343d659[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2cab66c3 (
    .a(al_281a7b5c),
    .b(al_4a463b38[28]),
    .c(al_794ac8f[9]),
    .o(al_e343d659[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f4f4898a (
    .a(al_281a7b5c),
    .b(al_4a463b38[29]),
    .c(al_794ac8f[10]),
    .o(al_e343d659[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9a7e1c26 (
    .a(al_281a7b5c),
    .b(al_4a463b38[30]),
    .c(al_794ac8f[11]),
    .o(al_e343d659[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3b425bcf (
    .a(al_281a7b5c),
    .b(al_4a463b38[31]),
    .c(al_794ac8f[12]),
    .o(al_e343d659[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e3632d2c (
    .a(al_281a7b5c),
    .b(al_4a463b38[32]),
    .c(al_794ac8f[13]),
    .o(al_e343d659[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fb39c8e (
    .a(al_281a7b5c),
    .b(al_4a463b38[33]),
    .c(al_794ac8f[14]),
    .o(al_e343d659[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_82fae575 (
    .a(al_281a7b5c),
    .b(al_4a463b38[34]),
    .c(al_794ac8f[15]),
    .o(al_e343d659[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e9f0092b (
    .a(al_281a7b5c),
    .b(al_4a463b38[35]),
    .c(al_794ac8f[16]),
    .o(al_e343d659[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7d5d1779 (
    .a(al_281a7b5c),
    .b(al_4a463b38[36]),
    .c(al_794ac8f[17]),
    .o(al_e343d659[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_58826389 (
    .a(al_281a7b5c),
    .b(al_4a463b38[37]),
    .c(al_794ac8f[18]),
    .o(al_e343d659[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_99b6585b (
    .a(al_281a7b5c),
    .b(al_4a463b38[38]),
    .c(al_794ac8f[19]),
    .o(al_e343d659[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5e7cc360 (
    .a(al_281a7b5c),
    .b(al_4a463b38[39]),
    .c(al_794ac8f[20]),
    .o(al_e343d659[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_75cea068 (
    .a(al_281a7b5c),
    .b(al_4a463b38[40]),
    .c(al_794ac8f[21]),
    .o(al_e343d659[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7b2a82d2 (
    .a(al_281a7b5c),
    .b(al_4a463b38[41]),
    .c(al_794ac8f[22]),
    .o(al_e343d659[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_31a194f6 (
    .a(al_281a7b5c),
    .b(al_4a463b38[42]),
    .c(al_794ac8f[23]),
    .o(al_e343d659[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_39d18360 (
    .a(al_281a7b5c),
    .b(al_4a463b38[43]),
    .c(al_794ac8f[24]),
    .o(al_e343d659[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8ed8773e (
    .a(al_281a7b5c),
    .b(al_4a463b38[44]),
    .c(al_794ac8f[25]),
    .o(al_e343d659[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8f84c1e4 (
    .a(al_281a7b5c),
    .b(al_4a463b38[45]),
    .c(al_794ac8f[26]),
    .o(al_e343d659[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_29dff70d (
    .a(al_281a7b5c),
    .b(al_4a463b38[46]),
    .c(al_794ac8f[27]),
    .o(al_e343d659[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bcebd93e (
    .a(al_281a7b5c),
    .b(al_4a463b38[47]),
    .c(al_794ac8f[28]),
    .o(al_e343d659[47]));
  AL_DFF_X al_3706542b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[0]));
  AL_DFF_X al_424c7aa8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[9]));
  AL_DFF_X al_8f40b476 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[10]));
  AL_DFF_X al_2169d00d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[11]));
  AL_DFF_X al_9844dccf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[12]));
  AL_DFF_X al_df363dd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[13]));
  AL_DFF_X al_cf4bbb4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[14]));
  AL_DFF_X al_a7dc38e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[15]));
  AL_DFF_X al_7d148c57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[16]));
  AL_DFF_X al_bae024b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[17]));
  AL_DFF_X al_c1db038f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[18]));
  AL_DFF_X al_aa74f95e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[1]));
  AL_DFF_X al_4111008a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[19]));
  AL_DFF_X al_7f0c94d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[20]));
  AL_DFF_X al_70d03947 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[21]));
  AL_DFF_X al_6c3c3b45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[22]));
  AL_DFF_X al_9bb53f2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[23]));
  AL_DFF_X al_b9d35153 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[24]));
  AL_DFF_X al_6ba2eeef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[25]));
  AL_DFF_X al_7988929a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[26]));
  AL_DFF_X al_f8c16e89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[27]));
  AL_DFF_X al_4a76c996 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[28]));
  AL_DFF_X al_5a5ea10b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[2]));
  AL_DFF_X al_1676afa7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[29]));
  AL_DFF_X al_7d462afe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[30]));
  AL_DFF_X al_f648c890 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[31]));
  AL_DFF_X al_25cd1c16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[32]));
  AL_DFF_X al_6ac62fdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[33]));
  AL_DFF_X al_45dbcb93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[34]));
  AL_DFF_X al_be48db53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[35]));
  AL_DFF_X al_dde5a999 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[36]));
  AL_DFF_X al_1a6e6fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[37]));
  AL_DFF_X al_3a42631d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[38]));
  AL_DFF_X al_b25bf98d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[3]));
  AL_DFF_X al_1e8d4d03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[39]));
  AL_DFF_X al_9564d8ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[40]));
  AL_DFF_X al_6c422925 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[41]));
  AL_DFF_X al_56b26b07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[42]));
  AL_DFF_X al_c351074b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[43]));
  AL_DFF_X al_bcb2a37f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[44]));
  AL_DFF_X al_5013ccdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[45]));
  AL_DFF_X al_33c59a9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[46]));
  AL_DFF_X al_76f35f60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e343d659[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[47]));
  AL_DFF_X al_3a8e0f73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[4]));
  AL_DFF_X al_537da286 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[5]));
  AL_DFF_X al_fa1bb280 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[6]));
  AL_DFF_X al_452c3206 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[7]));
  AL_DFF_X al_960cdcf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4a463b38[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32ba5b24[8]));
  AL_DFF_X al_4171056 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_281a7b5c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[0]));
  AL_DFF_X al_63662f1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[9]));
  AL_DFF_X al_2801daeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[10]));
  AL_DFF_X al_b3a95fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[11]));
  AL_DFF_X al_1a4efb99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[12]));
  AL_DFF_X al_484fd955 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[13]));
  AL_DFF_X al_6031043c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[14]));
  AL_DFF_X al_8ced292b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[15]));
  AL_DFF_X al_44a21302 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[16]));
  AL_DFF_X al_5dd60aea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[17]));
  AL_DFF_X al_8a087a89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[18]));
  AL_DFF_X al_de507879 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[1]));
  AL_DFF_X al_693a5ccf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[19]));
  AL_DFF_X al_7793239b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[20]));
  AL_DFF_X al_1a90e606 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[21]));
  AL_DFF_X al_b5f80121 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[22]));
  AL_DFF_X al_78f7e239 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[23]));
  AL_DFF_X al_df614077 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[24]));
  AL_DFF_X al_bb4bf59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[25]));
  AL_DFF_X al_9230206c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[26]));
  AL_DFF_X al_eeef28dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[27]));
  AL_DFF_X al_9baad285 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[28]));
  AL_DFF_X al_b9e3d82d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[2]));
  AL_DFF_X al_fe7e8899 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[3]));
  AL_DFF_X al_c1fa7bd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[4]));
  AL_DFF_X al_2440a64a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[5]));
  AL_DFF_X al_abfa7f75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[6]));
  AL_DFF_X al_55342b59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[7]));
  AL_DFF_X al_dfa4732e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7a3cd65[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bad3f013[8]));
  AL_DFF_X al_170fcbf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5db428bb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8d805738[0]));
  AL_DFF_X al_e361eef2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[17]));
  AL_DFF_X al_4286ca57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[18]));
  AL_DFF_X al_74c47359 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[19]));
  AL_DFF_X al_8eb5f6ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[20]));
  AL_DFF_X al_ba2921d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[21]));
  AL_DFF_X al_cc00a5c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[22]));
  AL_DFF_X al_3b59b20e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[23]));
  AL_DFF_X al_e5cafa87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[24]));
  AL_DFF_X al_25bde4af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[25]));
  AL_DFF_X al_a6dbc1a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[26]));
  AL_DFF_X al_173621c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[27]));
  AL_DFF_X al_3632ebdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[28]));
  AL_DFF_X al_5dba3c2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[29]));
  AL_DFF_X al_837e124 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[30]));
  AL_DFF_X al_e0d1c8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[31]));
  AL_DFF_X al_3264ffc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[32]));
  AL_DFF_X al_1583e93a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[33]));
  AL_DFF_X al_e27dbb04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[34]));
  AL_DFF_X al_5f5b4a6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[35]));
  AL_DFF_X al_3d2d5752 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[36]));
  AL_DFF_X al_b44dfd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[37]));
  AL_DFF_X al_9692fca6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[38]));
  AL_DFF_X al_78af6b5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[39]));
  AL_DFF_X al_84b7d5ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[40]));
  AL_DFF_X al_3c4e6ba0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[41]));
  AL_DFF_X al_3f129e4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[42]));
  AL_DFF_X al_98141092 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[43]));
  AL_DFF_X al_c22dcf19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[44]));
  AL_DFF_X al_1a803f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[45]));
  AL_DFF_X al_4b5a9919 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[46]));
  AL_DFF_X al_5b2a22bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[47]));
  AL_DFF_X al_74887d2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d1a07609[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_627988c3[48]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_9daf285a (
    .a(1'b0),
    .o({al_17661190,open_n116}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a4dc4972 (
    .a(al_32ba5b24[18]),
    .b(al_d1a07609[18]),
    .c(al_17661190),
    .o({al_ba73d945,al_af127331[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_467aebfe (
    .a(al_32ba5b24[19]),
    .b(al_d1a07609[19]),
    .c(al_ba73d945),
    .o({al_7e55c045,al_af127331[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_426a078b (
    .a(al_32ba5b24[20]),
    .b(al_d1a07609[20]),
    .c(al_7e55c045),
    .o({al_efd0595d,al_af127331[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f2fc5f83 (
    .a(al_32ba5b24[21]),
    .b(al_d1a07609[21]),
    .c(al_efd0595d),
    .o({al_83ddd85b,al_af127331[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6e89ffa (
    .a(al_32ba5b24[22]),
    .b(al_d1a07609[22]),
    .c(al_83ddd85b),
    .o({al_4697075e,al_af127331[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_73fdff75 (
    .a(al_32ba5b24[23]),
    .b(al_d1a07609[23]),
    .c(al_4697075e),
    .o({al_5ad7048f,al_af127331[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_48f94e0a (
    .a(al_32ba5b24[24]),
    .b(al_d1a07609[24]),
    .c(al_5ad7048f),
    .o({al_9071f0e5,al_af127331[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5c67348a (
    .a(al_32ba5b24[25]),
    .b(al_d1a07609[25]),
    .c(al_9071f0e5),
    .o({al_e5398263,al_af127331[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6baa6508 (
    .a(al_32ba5b24[26]),
    .b(al_d1a07609[26]),
    .c(al_e5398263),
    .o({al_b191d1e0,al_af127331[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9a6133dc (
    .a(al_32ba5b24[27]),
    .b(al_d1a07609[27]),
    .c(al_b191d1e0),
    .o({al_49a0e61d,al_af127331[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2f4d107e (
    .a(al_32ba5b24[28]),
    .b(al_d1a07609[28]),
    .c(al_49a0e61d),
    .o({al_86984010,al_af127331[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f16d2767 (
    .a(al_32ba5b24[29]),
    .b(al_d1a07609[29]),
    .c(al_86984010),
    .o({al_862cc7f8,al_af127331[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_689cf914 (
    .a(al_32ba5b24[30]),
    .b(al_d1a07609[30]),
    .c(al_862cc7f8),
    .o({al_b980f13c,al_af127331[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5ea99c28 (
    .a(al_32ba5b24[31]),
    .b(al_d1a07609[31]),
    .c(al_b980f13c),
    .o({al_db4a0b3b,al_af127331[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_92994423 (
    .a(al_32ba5b24[32]),
    .b(al_d1a07609[32]),
    .c(al_db4a0b3b),
    .o({al_b7c44457,al_af127331[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_316a3d63 (
    .a(al_32ba5b24[33]),
    .b(al_d1a07609[33]),
    .c(al_b7c44457),
    .o({al_c68c13d2,al_af127331[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bca987a0 (
    .a(al_32ba5b24[34]),
    .b(al_d1a07609[34]),
    .c(al_c68c13d2),
    .o({al_f144ba04,al_af127331[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b81943ed (
    .a(al_32ba5b24[35]),
    .b(al_d1a07609[35]),
    .c(al_f144ba04),
    .o({al_2e50ac1e,al_af127331[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a37b6bbc (
    .a(al_32ba5b24[36]),
    .b(al_d1a07609[36]),
    .c(al_2e50ac1e),
    .o({al_e418756e,al_af127331[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2f8afbe4 (
    .a(al_32ba5b24[37]),
    .b(al_d1a07609[37]),
    .c(al_e418756e),
    .o({al_8653cc11,al_af127331[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_24a2f970 (
    .a(al_32ba5b24[38]),
    .b(al_d1a07609[38]),
    .c(al_8653cc11),
    .o({al_fa5db848,al_af127331[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eda24a6b (
    .a(al_32ba5b24[39]),
    .b(al_d1a07609[39]),
    .c(al_fa5db848),
    .o({al_39ade860,al_af127331[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5f972b78 (
    .a(al_32ba5b24[40]),
    .b(al_d1a07609[40]),
    .c(al_39ade860),
    .o({al_7183147,al_af127331[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b4194b3b (
    .a(al_32ba5b24[41]),
    .b(al_d1a07609[41]),
    .c(al_7183147),
    .o({al_616fbe10,al_af127331[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_64d3b47c (
    .a(al_32ba5b24[42]),
    .b(al_d1a07609[42]),
    .c(al_616fbe10),
    .o({al_47d76c66,al_af127331[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4f0d89be (
    .a(al_32ba5b24[43]),
    .b(al_d1a07609[43]),
    .c(al_47d76c66),
    .o({al_ebfbc5f1,al_af127331[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5379bc02 (
    .a(al_32ba5b24[44]),
    .b(al_d1a07609[44]),
    .c(al_ebfbc5f1),
    .o({al_3f596b4e,al_af127331[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f6a9933 (
    .a(al_32ba5b24[45]),
    .b(al_d1a07609[45]),
    .c(al_3f596b4e),
    .o({al_4b8b49e0,al_af127331[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cd86da99 (
    .a(al_32ba5b24[46]),
    .b(al_d1a07609[46]),
    .c(al_4b8b49e0),
    .o({al_608458c0,al_af127331[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d908b61c (
    .a(al_32ba5b24[47]),
    .b(al_d1a07609[47]),
    .c(al_608458c0),
    .o({al_14b22db9,al_af127331[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bdbe86b2 (
    .c(al_14b22db9),
    .o({open_n119,al_af127331[30]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_239f1f05 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[18]),
    .c(al_af127331[0]),
    .o(al_14165a56[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c07aa2d5 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[19]),
    .c(al_af127331[1]),
    .o(al_14165a56[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f445c83 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[20]),
    .c(al_af127331[2]),
    .o(al_14165a56[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_caf5d5cc (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[21]),
    .c(al_af127331[3]),
    .o(al_14165a56[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1769f616 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[22]),
    .c(al_af127331[4]),
    .o(al_14165a56[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7c92af4d (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[23]),
    .c(al_af127331[5]),
    .o(al_14165a56[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8a1fbdd (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[24]),
    .c(al_af127331[6]),
    .o(al_14165a56[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e8a834a0 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[25]),
    .c(al_af127331[7]),
    .o(al_14165a56[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_50cbb86b (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[26]),
    .c(al_af127331[8]),
    .o(al_14165a56[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f80656e (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[27]),
    .c(al_af127331[9]),
    .o(al_14165a56[27]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_e98bab02 (
    .a(al_d1a07609[48]),
    .b(al_d1a07609[49]),
    .c(al_af127331[30]),
    .o(al_f04c5c1a));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c6e86ff4 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[28]),
    .c(al_af127331[10]),
    .o(al_14165a56[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6080847d (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[29]),
    .c(al_af127331[11]),
    .o(al_14165a56[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4209a834 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[30]),
    .c(al_af127331[12]),
    .o(al_14165a56[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ddfa8cc3 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[31]),
    .c(al_af127331[13]),
    .o(al_14165a56[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2979ea73 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[32]),
    .c(al_af127331[14]),
    .o(al_14165a56[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_84acf2d1 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[33]),
    .c(al_af127331[15]),
    .o(al_14165a56[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fbf13339 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[34]),
    .c(al_af127331[16]),
    .o(al_14165a56[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_45e39180 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[35]),
    .c(al_af127331[17]),
    .o(al_14165a56[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_12ddc882 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[36]),
    .c(al_af127331[18]),
    .o(al_14165a56[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6b752df7 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[37]),
    .c(al_af127331[19]),
    .o(al_14165a56[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dc05b54b (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[38]),
    .c(al_af127331[20]),
    .o(al_14165a56[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_49fa2171 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[39]),
    .c(al_af127331[21]),
    .o(al_14165a56[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_606a38d7 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[40]),
    .c(al_af127331[22]),
    .o(al_14165a56[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_fe3c95ae (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[41]),
    .c(al_af127331[23]),
    .o(al_14165a56[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2c8c04a1 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[42]),
    .c(al_af127331[24]),
    .o(al_14165a56[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5fd78972 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[43]),
    .c(al_af127331[25]),
    .o(al_14165a56[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ad20de2e (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[44]),
    .c(al_af127331[26]),
    .o(al_14165a56[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_51a2d171 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[45]),
    .c(al_af127331[27]),
    .o(al_14165a56[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_97e32dfc (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[46]),
    .c(al_af127331[28]),
    .o(al_14165a56[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_332b94b8 (
    .a(al_f04c5c1a),
    .b(al_32ba5b24[47]),
    .c(al_af127331[29]),
    .o(al_14165a56[47]));
  AL_DFF_X al_cd94e03a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[0]));
  AL_DFF_X al_21d805c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[9]));
  AL_DFF_X al_1379d2d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[10]));
  AL_DFF_X al_970129bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[11]));
  AL_DFF_X al_aae212d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[12]));
  AL_DFF_X al_2b722404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[13]));
  AL_DFF_X al_411274a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[14]));
  AL_DFF_X al_712f88fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[15]));
  AL_DFF_X al_e79edad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[16]));
  AL_DFF_X al_f8048dec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[17]));
  AL_DFF_X al_f77418d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[18]));
  AL_DFF_X al_25a3e905 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[1]));
  AL_DFF_X al_b8a8cc84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[19]));
  AL_DFF_X al_b84551fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[20]));
  AL_DFF_X al_71cff4c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[21]));
  AL_DFF_X al_4a80d1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[22]));
  AL_DFF_X al_e307e7dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[23]));
  AL_DFF_X al_11e212dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[24]));
  AL_DFF_X al_5daade08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[25]));
  AL_DFF_X al_2a002d46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[26]));
  AL_DFF_X al_6c6787c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[27]));
  AL_DFF_X al_a895e22d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[28]));
  AL_DFF_X al_b2c4958b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[2]));
  AL_DFF_X al_46615397 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[29]));
  AL_DFF_X al_99e988bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[30]));
  AL_DFF_X al_a0c8f676 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[31]));
  AL_DFF_X al_b100cdf2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[32]));
  AL_DFF_X al_fa94be25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[33]));
  AL_DFF_X al_e6048909 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[34]));
  AL_DFF_X al_443733d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[35]));
  AL_DFF_X al_269cba6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[36]));
  AL_DFF_X al_f901bc6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[37]));
  AL_DFF_X al_ac536b83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[38]));
  AL_DFF_X al_f743ac7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[3]));
  AL_DFF_X al_ce2dbf32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[39]));
  AL_DFF_X al_3a03023a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[40]));
  AL_DFF_X al_d5f70bff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[41]));
  AL_DFF_X al_69f6cf6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[42]));
  AL_DFF_X al_cadb88c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[43]));
  AL_DFF_X al_a8421eed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[44]));
  AL_DFF_X al_a3ed9ff9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[45]));
  AL_DFF_X al_39219bdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[46]));
  AL_DFF_X al_d59d1ee5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_14165a56[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[47]));
  AL_DFF_X al_3d7a7a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[4]));
  AL_DFF_X al_f6b8df91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[5]));
  AL_DFF_X al_39dce3d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[6]));
  AL_DFF_X al_4dc1291b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[7]));
  AL_DFF_X al_5feccb95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32ba5b24[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_690b21a4[8]));
  AL_DFF_X al_2b7f0f1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f04c5c1a),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[0]));
  AL_DFF_X al_fa44b1ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[9]));
  AL_DFF_X al_8fd83b53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[10]));
  AL_DFF_X al_4df80905 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[11]));
  AL_DFF_X al_92fe1c30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[12]));
  AL_DFF_X al_5edcab9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[13]));
  AL_DFF_X al_799920cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[14]));
  AL_DFF_X al_55783b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[15]));
  AL_DFF_X al_a24db40c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[16]));
  AL_DFF_X al_39a12728 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[17]));
  AL_DFF_X al_1a3a20ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[18]));
  AL_DFF_X al_66b87332 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[1]));
  AL_DFF_X al_a5aedaef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[19]));
  AL_DFF_X al_f2a0ee0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[20]));
  AL_DFF_X al_15cc2784 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[21]));
  AL_DFF_X al_d915116f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[22]));
  AL_DFF_X al_5d58cedd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[23]));
  AL_DFF_X al_653f755b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[24]));
  AL_DFF_X al_d7945c2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[25]));
  AL_DFF_X al_89bc922 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[26]));
  AL_DFF_X al_d877dd06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[27]));
  AL_DFF_X al_1bda18dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[28]));
  AL_DFF_X al_a24676df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[2]));
  AL_DFF_X al_d80f064e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[29]));
  AL_DFF_X al_f381c8a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[3]));
  AL_DFF_X al_1072b16c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[4]));
  AL_DFF_X al_8bacdf39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[5]));
  AL_DFF_X al_4592713f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[6]));
  AL_DFF_X al_13a820c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[7]));
  AL_DFF_X al_414b0833 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bad3f013[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d67405f[8]));
  AL_DFF_X al_3d9f134d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_67f5b0b3[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44882eca[0]));
  AL_DFF_X al_74beed6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[44]));
  AL_DFF_X al_a0f807ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[45]));
  AL_DFF_X al_e3354ee4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[46]));
  AL_DFF_X al_7a949f96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[47]));
  AL_DFF_X al_80460a73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[48]));
  AL_DFF_X al_8ecdcc30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[49]));
  AL_DFF_X al_5b76812a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[50]));
  AL_DFF_X al_ff2e216a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[51]));
  AL_DFF_X al_906a1d70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[52]));
  AL_DFF_X al_60d2d1e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[53]));
  AL_DFF_X al_b2cd76bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[54]));
  AL_DFF_X al_48280716 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[55]));
  AL_DFF_X al_5151c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[56]));
  AL_DFF_X al_a363277b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[57]));
  AL_DFF_X al_9ed07d73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[58]));
  AL_DFF_X al_77f6c9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[59]));
  AL_DFF_X al_4ec1f27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[60]));
  AL_DFF_X al_56da25a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[61]));
  AL_DFF_X al_6a98fec2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[62]));
  AL_DFF_X al_d2872c90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[63]));
  AL_DFF_X al_d0c04a35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[64]));
  AL_DFF_X al_821f83db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[65]));
  AL_DFF_X al_8530ed8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[66]));
  AL_DFF_X al_5916251 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[67]));
  AL_DFF_X al_884bfaac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[68]));
  AL_DFF_X al_c678633d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[69]));
  AL_DFF_X al_cee3823a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[70]));
  AL_DFF_X al_9c8b8073 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[71]));
  AL_DFF_X al_190a94de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[72]));
  AL_DFF_X al_1f730d97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[73]));
  AL_DFF_X al_1350832e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[74]));
  AL_DFF_X al_fde06bc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6a637a32[76]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b052c226[75]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_ea578487 (
    .a(al_b34ec3bf),
    .b(al_2aef1337),
    .o(al_ffbd9e7e));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    al_ea48af86 (
    .a(al_6a637a32[45]),
    .b(al_3d0cfeb4[45]),
    .o(al_b33cc591));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_d0b122df (
    .a(al_6a637a32[48]),
    .b(al_6a637a32[49]),
    .o(al_1c1f1cb1));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_c4a62743 (
    .a(al_6a637a32[56]),
    .b(al_6a637a32[57]),
    .c(al_6a637a32[58]),
    .d(al_6a637a32[59]),
    .e(al_6a637a32[60]),
    .f(al_6a637a32[61]),
    .o(al_55f734a7));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_2db3287f (
    .a(al_6a637a32[50]),
    .b(al_6a637a32[51]),
    .c(al_6a637a32[52]),
    .d(al_6a637a32[53]),
    .e(al_6a637a32[54]),
    .f(al_6a637a32[55]),
    .o(al_51e8603));
  AL_MAP_LUT6 #(
    .EQN("(F*E*D*C*B*A)"),
    .INIT(64'h8000000000000000))
    al_656e51a7 (
    .a(al_eb58c5cb),
    .b(al_95542881),
    .c(al_8b31dee3),
    .d(al_1c1f1cb1),
    .e(al_55f734a7),
    .f(al_51e8603),
    .o(al_2aef1337));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*B*~A))"),
    .INIT(16'hbf40))
    al_f4c8f342 (
    .a(al_b34ec3bf),
    .b(al_2aef1337),
    .c(al_6a637a32[45]),
    .d(al_3d0cfeb4[45]),
    .o(al_a9b28455[45]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*B*C*D*E)"),
    .INIT(32'h80e0f8fe))
    al_16ba429c (
    .a(al_b33cc591),
    .b(al_6a637a32[46]),
    .c(al_6a637a32[47]),
    .d(al_3d0cfeb4[46]),
    .e(al_3d0cfeb4[47]),
    .o(al_b34ec3bf));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_e3dccc08 (
    .a(al_6a637a32[70]),
    .b(al_6a637a32[71]),
    .c(al_6a637a32[72]),
    .d(al_6a637a32[73]),
    .e(al_6a637a32[74]),
    .f(al_6a637a32[75]),
    .o(al_eb58c5cb));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_eac6388a (
    .a(al_6a637a32[64]),
    .b(al_6a637a32[65]),
    .c(al_6a637a32[66]),
    .d(al_6a637a32[67]),
    .e(al_6a637a32[68]),
    .f(al_6a637a32[69]),
    .o(al_95542881));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_2a183cbf (
    .a(al_6a637a32[62]),
    .b(al_6a637a32[63]),
    .c(al_6a637a32[76]),
    .o(al_8b31dee3));
  AL_MAP_LUT5 #(
    .EQN("(D*C*B*(E@A))"),
    .INIT(32'h40008000))
    al_7b8bba2d (
    .a(al_b33cc591),
    .b(al_eb58c5cb),
    .c(al_95542881),
    .d(al_8b31dee3),
    .e(al_6a637a32[46]),
    .o(al_6b3dc9d));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_749f75bc (
    .a(al_b34ec3bf),
    .b(al_6b3dc9d),
    .c(al_1c1f1cb1),
    .d(al_55f734a7),
    .e(al_51e8603),
    .f(al_3d0cfeb4[46]),
    .o(al_a9b28455[46]));
  AL_MAP_LUT6 #(
    .EQN("(F*~(A*~(D@(~(B)*~(C)*~(E)+~(B)*~(C)*E+B*~(C)*E+~(B)*C*E))))"),
    .INIT(64'hd57ffd5700000000))
    al_91984e56 (
    .a(al_2aef1337),
    .b(al_b33cc591),
    .c(al_6a637a32[46]),
    .d(al_6a637a32[47]),
    .e(al_3d0cfeb4[46]),
    .f(al_3d0cfeb4[47]),
    .o(al_a9b28455[47]));
  AL_DFF_X al_71778710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[0]));
  AL_DFF_X al_5d309d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[9]));
  AL_DFF_X al_2237bf28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[10]));
  AL_DFF_X al_fc30d591 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[11]));
  AL_DFF_X al_99f6132d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[12]));
  AL_DFF_X al_37ddf104 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[13]));
  AL_DFF_X al_4d42dc67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[14]));
  AL_DFF_X al_ad449795 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[15]));
  AL_DFF_X al_8bc31585 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[16]));
  AL_DFF_X al_7b42e7c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[17]));
  AL_DFF_X al_d5d15018 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[18]));
  AL_DFF_X al_a5449fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[1]));
  AL_DFF_X al_c7a7ddd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[19]));
  AL_DFF_X al_c2844f7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[20]));
  AL_DFF_X al_2bebe6ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[21]));
  AL_DFF_X al_9baa590c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[22]));
  AL_DFF_X al_4de1ff33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[23]));
  AL_DFF_X al_7db2c016 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[24]));
  AL_DFF_X al_58e14091 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[25]));
  AL_DFF_X al_42465b64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[26]));
  AL_DFF_X al_836ed255 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[27]));
  AL_DFF_X al_c587b35c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[28]));
  AL_DFF_X al_9376a561 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[2]));
  AL_DFF_X al_48136e64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[29]));
  AL_DFF_X al_3579d0cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[30]));
  AL_DFF_X al_31afc303 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[31]));
  AL_DFF_X al_9556f8cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[32]));
  AL_DFF_X al_78e67288 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[33]));
  AL_DFF_X al_56c67f97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[34]));
  AL_DFF_X al_ba9d3c81 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[35]));
  AL_DFF_X al_9726ff2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[36]));
  AL_DFF_X al_e52fe31d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[37]));
  AL_DFF_X al_caa2f87a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[38]));
  AL_DFF_X al_c44982f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[3]));
  AL_DFF_X al_13852169 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[39]));
  AL_DFF_X al_d1b62590 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[40]));
  AL_DFF_X al_711cb688 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[41]));
  AL_DFF_X al_7c1bca5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[42]));
  AL_DFF_X al_d9e3d02c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[43]));
  AL_DFF_X al_1f726616 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[44]));
  AL_DFF_X al_6cf6c769 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9b28455[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[45]));
  AL_DFF_X al_a0b6f109 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9b28455[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[46]));
  AL_DFF_X al_e92808b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a9b28455[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[47]));
  AL_DFF_X al_fe0fb942 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[4]));
  AL_DFF_X al_227282d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[5]));
  AL_DFF_X al_8efbe81b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[6]));
  AL_DFF_X al_6036d0ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[7]));
  AL_DFF_X al_5dd53115 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3d0cfeb4[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_592f1b09[8]));
  AL_DFF_X al_969f6ae5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ffbd9e7e),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b18b7cbb[0]));
  AL_DFF_X al_b6f7f69c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b54c1014[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b18b7cbb[1]));
  AL_DFF_X al_178b777f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b54c1014[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b18b7cbb[2]));
  AL_DFF_X al_cd0a560a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8d805738[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_74993dd2[0]));
  AL_DFF_X al_eafb9dcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[16]));
  AL_DFF_X al_26a6750c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[17]));
  AL_DFF_X al_48d28b1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[18]));
  AL_DFF_X al_342d2606 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[19]));
  AL_DFF_X al_4db46a23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[20]));
  AL_DFF_X al_eee162b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[21]));
  AL_DFF_X al_a8e62efc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[22]));
  AL_DFF_X al_f46b98f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[23]));
  AL_DFF_X al_d3385f6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[24]));
  AL_DFF_X al_b329a79c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[25]));
  AL_DFF_X al_f081e8c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[26]));
  AL_DFF_X al_e661b646 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[27]));
  AL_DFF_X al_c4e3d6b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[28]));
  AL_DFF_X al_b6a563cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[29]));
  AL_DFF_X al_9d6f264d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[30]));
  AL_DFF_X al_4e656419 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[31]));
  AL_DFF_X al_e6cf4b9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[32]));
  AL_DFF_X al_3b66a355 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[33]));
  AL_DFF_X al_56edb17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[34]));
  AL_DFF_X al_75086750 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[35]));
  AL_DFF_X al_17d5777 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[36]));
  AL_DFF_X al_7eea3b06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[37]));
  AL_DFF_X al_f29b6392 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[38]));
  AL_DFF_X al_4027e7ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[39]));
  AL_DFF_X al_7aca0448 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[40]));
  AL_DFF_X al_7fbb5d42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[41]));
  AL_DFF_X al_b0ebaec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[42]));
  AL_DFF_X al_fec57970 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[43]));
  AL_DFF_X al_bd95a5d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[44]));
  AL_DFF_X al_2a431e30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[45]));
  AL_DFF_X al_437a51d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[46]));
  AL_DFF_X al_b24955b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_627988c3[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5e9c08d[47]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_7a6c4e19 (
    .a(1'b0),
    .o({al_a3fc3ebc,open_n122}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b3131dc6 (
    .a(al_690b21a4[17]),
    .b(al_627988c3[17]),
    .c(al_a3fc3ebc),
    .o({al_5cdd85d5,al_2c47200f[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1480afec (
    .a(al_690b21a4[18]),
    .b(al_627988c3[18]),
    .c(al_5cdd85d5),
    .o({al_1add508,al_2c47200f[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67773c4e (
    .a(al_690b21a4[19]),
    .b(al_627988c3[19]),
    .c(al_1add508),
    .o({al_5a84d22c,al_2c47200f[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_daee945f (
    .a(al_690b21a4[20]),
    .b(al_627988c3[20]),
    .c(al_5a84d22c),
    .o({al_cf720ce3,al_2c47200f[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bf9fcca (
    .a(al_690b21a4[21]),
    .b(al_627988c3[21]),
    .c(al_cf720ce3),
    .o({al_656d5c84,al_2c47200f[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d75f392d (
    .a(al_690b21a4[22]),
    .b(al_627988c3[22]),
    .c(al_656d5c84),
    .o({al_de32c090,al_2c47200f[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3484982 (
    .a(al_690b21a4[23]),
    .b(al_627988c3[23]),
    .c(al_de32c090),
    .o({al_f42fa6ce,al_2c47200f[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67a80a6d (
    .a(al_690b21a4[24]),
    .b(al_627988c3[24]),
    .c(al_f42fa6ce),
    .o({al_b6af5571,al_2c47200f[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fa781ea6 (
    .a(al_690b21a4[25]),
    .b(al_627988c3[25]),
    .c(al_b6af5571),
    .o({al_c2ee5e5b,al_2c47200f[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2ee5b555 (
    .a(al_690b21a4[26]),
    .b(al_627988c3[26]),
    .c(al_c2ee5e5b),
    .o({al_43f00cc1,al_2c47200f[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b85ee9a0 (
    .a(al_690b21a4[27]),
    .b(al_627988c3[27]),
    .c(al_43f00cc1),
    .o({al_a541ec8a,al_2c47200f[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_da58d88e (
    .a(al_690b21a4[28]),
    .b(al_627988c3[28]),
    .c(al_a541ec8a),
    .o({al_74501eb3,al_2c47200f[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3373ae9a (
    .a(al_690b21a4[29]),
    .b(al_627988c3[29]),
    .c(al_74501eb3),
    .o({al_ffc5f376,al_2c47200f[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5d90a9e8 (
    .a(al_690b21a4[30]),
    .b(al_627988c3[30]),
    .c(al_ffc5f376),
    .o({al_d3b64099,al_2c47200f[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ab7e3864 (
    .a(al_690b21a4[31]),
    .b(al_627988c3[31]),
    .c(al_d3b64099),
    .o({al_9abafd70,al_2c47200f[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_16e73e4c (
    .a(al_690b21a4[32]),
    .b(al_627988c3[32]),
    .c(al_9abafd70),
    .o({al_8225507c,al_2c47200f[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4b24d558 (
    .a(al_690b21a4[33]),
    .b(al_627988c3[33]),
    .c(al_8225507c),
    .o({al_ff92482,al_2c47200f[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_420d2cce (
    .a(al_690b21a4[34]),
    .b(al_627988c3[34]),
    .c(al_ff92482),
    .o({al_2e13f976,al_2c47200f[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f33da7d9 (
    .a(al_690b21a4[35]),
    .b(al_627988c3[35]),
    .c(al_2e13f976),
    .o({al_bd65eabf,al_2c47200f[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_55c9af34 (
    .a(al_690b21a4[36]),
    .b(al_627988c3[36]),
    .c(al_bd65eabf),
    .o({al_ede5673b,al_2c47200f[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_78cae2e8 (
    .a(al_690b21a4[37]),
    .b(al_627988c3[37]),
    .c(al_ede5673b),
    .o({al_70a9c221,al_2c47200f[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9aad8383 (
    .a(al_690b21a4[38]),
    .b(al_627988c3[38]),
    .c(al_70a9c221),
    .o({al_532cc9a8,al_2c47200f[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ac55b8c1 (
    .a(al_690b21a4[39]),
    .b(al_627988c3[39]),
    .c(al_532cc9a8),
    .o({al_ea82bb3a,al_2c47200f[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7d5c9c15 (
    .a(al_690b21a4[40]),
    .b(al_627988c3[40]),
    .c(al_ea82bb3a),
    .o({al_d637b77b,al_2c47200f[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_963ff519 (
    .a(al_690b21a4[41]),
    .b(al_627988c3[41]),
    .c(al_d637b77b),
    .o({al_2e7f5ba5,al_2c47200f[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_79f79d19 (
    .a(al_690b21a4[42]),
    .b(al_627988c3[42]),
    .c(al_2e7f5ba5),
    .o({al_93b7a367,al_2c47200f[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cfb625d (
    .a(al_690b21a4[43]),
    .b(al_627988c3[43]),
    .c(al_93b7a367),
    .o({al_3d8d5fa3,al_2c47200f[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f4fca905 (
    .a(al_690b21a4[44]),
    .b(al_627988c3[44]),
    .c(al_3d8d5fa3),
    .o({al_294cc864,al_2c47200f[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_627ffead (
    .a(al_690b21a4[45]),
    .b(al_627988c3[45]),
    .c(al_294cc864),
    .o({al_3220468,al_2c47200f[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d24c753b (
    .a(al_690b21a4[46]),
    .b(al_627988c3[46]),
    .c(al_3220468),
    .o({al_b1e53313,al_2c47200f[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e8194b00 (
    .a(al_690b21a4[47]),
    .b(al_627988c3[47]),
    .c(al_b1e53313),
    .o({al_e4e8fccd,al_2c47200f[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7be0f383 (
    .c(al_e4e8fccd),
    .o({open_n125,al_2c47200f[31]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_971e1476 (
    .a(al_d45bda05),
    .b(al_690b21a4[17]),
    .c(al_2c47200f[0]),
    .o(al_3ccb3a4f[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_912b0dd0 (
    .a(al_d45bda05),
    .b(al_690b21a4[18]),
    .c(al_2c47200f[1]),
    .o(al_3ccb3a4f[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_da7f19aa (
    .a(al_d45bda05),
    .b(al_690b21a4[19]),
    .c(al_2c47200f[2]),
    .o(al_3ccb3a4f[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_329f04d4 (
    .a(al_d45bda05),
    .b(al_690b21a4[20]),
    .c(al_2c47200f[3]),
    .o(al_3ccb3a4f[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_38fb5244 (
    .a(al_d45bda05),
    .b(al_690b21a4[21]),
    .c(al_2c47200f[4]),
    .o(al_3ccb3a4f[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b77668a5 (
    .a(al_d45bda05),
    .b(al_690b21a4[22]),
    .c(al_2c47200f[5]),
    .o(al_3ccb3a4f[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_b0a229ca (
    .a(al_d45bda05),
    .b(al_690b21a4[23]),
    .c(al_2c47200f[6]),
    .o(al_3ccb3a4f[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f62d7f63 (
    .a(al_d45bda05),
    .b(al_690b21a4[24]),
    .c(al_2c47200f[7]),
    .o(al_3ccb3a4f[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7583c301 (
    .a(al_d45bda05),
    .b(al_690b21a4[25]),
    .c(al_2c47200f[8]),
    .o(al_3ccb3a4f[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_505a1d48 (
    .a(al_d45bda05),
    .b(al_690b21a4[26]),
    .c(al_2c47200f[9]),
    .o(al_3ccb3a4f[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_bd67a4d5 (
    .a(al_d45bda05),
    .b(al_690b21a4[27]),
    .c(al_2c47200f[10]),
    .o(al_3ccb3a4f[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9d2c0b95 (
    .a(al_d45bda05),
    .b(al_690b21a4[28]),
    .c(al_2c47200f[11]),
    .o(al_3ccb3a4f[28]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    al_667996f6 (
    .a(al_627988c3[48]),
    .b(al_2c47200f[31]),
    .o(al_d45bda05));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8a73c4a5 (
    .a(al_d45bda05),
    .b(al_690b21a4[29]),
    .c(al_2c47200f[12]),
    .o(al_3ccb3a4f[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9e4c789e (
    .a(al_d45bda05),
    .b(al_690b21a4[30]),
    .c(al_2c47200f[13]),
    .o(al_3ccb3a4f[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f4400b70 (
    .a(al_d45bda05),
    .b(al_690b21a4[31]),
    .c(al_2c47200f[14]),
    .o(al_3ccb3a4f[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_37101e2d (
    .a(al_d45bda05),
    .b(al_690b21a4[32]),
    .c(al_2c47200f[15]),
    .o(al_3ccb3a4f[32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6a6e7ead (
    .a(al_d45bda05),
    .b(al_690b21a4[33]),
    .c(al_2c47200f[16]),
    .o(al_3ccb3a4f[33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a1bf94f8 (
    .a(al_d45bda05),
    .b(al_690b21a4[34]),
    .c(al_2c47200f[17]),
    .o(al_3ccb3a4f[34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cde71bbf (
    .a(al_d45bda05),
    .b(al_690b21a4[35]),
    .c(al_2c47200f[18]),
    .o(al_3ccb3a4f[35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2952e50b (
    .a(al_d45bda05),
    .b(al_690b21a4[36]),
    .c(al_2c47200f[19]),
    .o(al_3ccb3a4f[36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6dc38519 (
    .a(al_d45bda05),
    .b(al_690b21a4[37]),
    .c(al_2c47200f[20]),
    .o(al_3ccb3a4f[37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_edc56307 (
    .a(al_d45bda05),
    .b(al_690b21a4[38]),
    .c(al_2c47200f[21]),
    .o(al_3ccb3a4f[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a2a9298f (
    .a(al_d45bda05),
    .b(al_690b21a4[39]),
    .c(al_2c47200f[22]),
    .o(al_3ccb3a4f[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_88d55180 (
    .a(al_d45bda05),
    .b(al_690b21a4[40]),
    .c(al_2c47200f[23]),
    .o(al_3ccb3a4f[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ef2eb719 (
    .a(al_d45bda05),
    .b(al_690b21a4[41]),
    .c(al_2c47200f[24]),
    .o(al_3ccb3a4f[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dfb02a1 (
    .a(al_d45bda05),
    .b(al_690b21a4[42]),
    .c(al_2c47200f[25]),
    .o(al_3ccb3a4f[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_478e7894 (
    .a(al_d45bda05),
    .b(al_690b21a4[43]),
    .c(al_2c47200f[26]),
    .o(al_3ccb3a4f[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_dfee17f (
    .a(al_d45bda05),
    .b(al_690b21a4[44]),
    .c(al_2c47200f[27]),
    .o(al_3ccb3a4f[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3b86b9c6 (
    .a(al_d45bda05),
    .b(al_690b21a4[45]),
    .c(al_2c47200f[28]),
    .o(al_3ccb3a4f[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_124ee46a (
    .a(al_d45bda05),
    .b(al_690b21a4[46]),
    .c(al_2c47200f[29]),
    .o(al_3ccb3a4f[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_176a355f (
    .a(al_d45bda05),
    .b(al_690b21a4[47]),
    .c(al_2c47200f[30]),
    .o(al_3ccb3a4f[47]));
  AL_DFF_X al_dbc55c6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[0]));
  AL_DFF_X al_6315348b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[9]));
  AL_DFF_X al_b1dcdbe5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[10]));
  AL_DFF_X al_103e6c20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[11]));
  AL_DFF_X al_f64710e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[12]));
  AL_DFF_X al_b17c4977 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[13]));
  AL_DFF_X al_13ddc4ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[14]));
  AL_DFF_X al_e35eb15f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[15]));
  AL_DFF_X al_363378e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[16]));
  AL_DFF_X al_61b51f28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[17]));
  AL_DFF_X al_cd23054a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[18]));
  AL_DFF_X al_1e012f14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[1]));
  AL_DFF_X al_da7e98e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[19]));
  AL_DFF_X al_964c75c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[20]));
  AL_DFF_X al_9f300511 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[21]));
  AL_DFF_X al_ce28f8a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[22]));
  AL_DFF_X al_58eeab7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[23]));
  AL_DFF_X al_5b8bb64e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[24]));
  AL_DFF_X al_734fec53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[25]));
  AL_DFF_X al_ac3a9476 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[26]));
  AL_DFF_X al_68a2e2f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[27]));
  AL_DFF_X al_a71b29c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[28]));
  AL_DFF_X al_b68b98c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[2]));
  AL_DFF_X al_7d4f7cbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[29]));
  AL_DFF_X al_ab19bbcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[30]));
  AL_DFF_X al_75fd8aef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[31]));
  AL_DFF_X al_aabf597d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[32]));
  AL_DFF_X al_b93cd3a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[33]));
  AL_DFF_X al_466cf3ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[34]));
  AL_DFF_X al_8926e788 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[35]));
  AL_DFF_X al_a44273c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[36]));
  AL_DFF_X al_3ea2b01b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[37]));
  AL_DFF_X al_7b5e124a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[38]));
  AL_DFF_X al_8f8b01c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[3]));
  AL_DFF_X al_c2928501 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[39]));
  AL_DFF_X al_b8cf56cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[40]));
  AL_DFF_X al_e611c560 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[41]));
  AL_DFF_X al_9dcf102a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[42]));
  AL_DFF_X al_6b77b02a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[43]));
  AL_DFF_X al_4d411626 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[44]));
  AL_DFF_X al_15401a1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[45]));
  AL_DFF_X al_89dba604 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[46]));
  AL_DFF_X al_bbf27e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3ccb3a4f[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[47]));
  AL_DFF_X al_b5c88d4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[4]));
  AL_DFF_X al_879a5839 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[5]));
  AL_DFF_X al_da143ebc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[6]));
  AL_DFF_X al_74f0518d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[7]));
  AL_DFF_X al_a7a1f460 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_690b21a4[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_57dc9b0c[8]));
  AL_DFF_X al_f955fe4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d45bda05),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[0]));
  AL_DFF_X al_3ee3e06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[9]));
  AL_DFF_X al_71c6a847 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[10]));
  AL_DFF_X al_7cd172b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[11]));
  AL_DFF_X al_195340c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[12]));
  AL_DFF_X al_20f4f161 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[13]));
  AL_DFF_X al_e8994277 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[14]));
  AL_DFF_X al_a46a052 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[15]));
  AL_DFF_X al_46fba005 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[16]));
  AL_DFF_X al_e05ab842 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[17]));
  AL_DFF_X al_7f2861d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[18]));
  AL_DFF_X al_e68f450b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[1]));
  AL_DFF_X al_1a3e195c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[19]));
  AL_DFF_X al_fab597f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[20]));
  AL_DFF_X al_557744e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[21]));
  AL_DFF_X al_1b7a0522 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[22]));
  AL_DFF_X al_ab42c93a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[23]));
  AL_DFF_X al_a1bce4af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[24]));
  AL_DFF_X al_5400cf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[25]));
  AL_DFF_X al_f9a1ef25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[26]));
  AL_DFF_X al_56fd5621 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[27]));
  AL_DFF_X al_7a92a39c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[28]));
  AL_DFF_X al_1bc05d54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[2]));
  AL_DFF_X al_c410cc5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[29]));
  AL_DFF_X al_492fbcdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[30]));
  AL_DFF_X al_29a7ae9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[3]));
  AL_DFF_X al_212dc787 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[4]));
  AL_DFF_X al_187bfcf8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[5]));
  AL_DFF_X al_5973db71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[6]));
  AL_DFF_X al_a4db90d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[7]));
  AL_DFF_X al_64019223 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9d67405f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b40233aa[8]));
  AL_DFF_X al_752f9ec3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_74993dd2[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2e2a074f[0]));
  AL_DFF_X al_4461e0fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[15]));
  AL_DFF_X al_abeee547 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[16]));
  AL_DFF_X al_3b36ffd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[17]));
  AL_DFF_X al_c20bb553 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[18]));
  AL_DFF_X al_72667039 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[19]));
  AL_DFF_X al_da8faf9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[20]));
  AL_DFF_X al_88848090 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[21]));
  AL_DFF_X al_2b82e15a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[22]));
  AL_DFF_X al_1e8c6831 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[23]));
  AL_DFF_X al_fd525f72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[24]));
  AL_DFF_X al_280a9005 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[25]));
  AL_DFF_X al_3dd9196b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[26]));
  AL_DFF_X al_aec62f54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[27]));
  AL_DFF_X al_cca094fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[28]));
  AL_DFF_X al_dd149ab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[29]));
  AL_DFF_X al_161e82da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[30]));
  AL_DFF_X al_b37acecc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[31]));
  AL_DFF_X al_5e0d0334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[32]));
  AL_DFF_X al_5a6d9d83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[33]));
  AL_DFF_X al_616b1c07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[34]));
  AL_DFF_X al_3c9eedeb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[35]));
  AL_DFF_X al_d2ae0493 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[36]));
  AL_DFF_X al_6ddc179c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[37]));
  AL_DFF_X al_40ba97a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[38]));
  AL_DFF_X al_a81b39aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[39]));
  AL_DFF_X al_a83be6b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[40]));
  AL_DFF_X al_169c1823 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[41]));
  AL_DFF_X al_38a5bf64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[42]));
  AL_DFF_X al_9aeb3aec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[43]));
  AL_DFF_X al_27c86cfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[44]));
  AL_DFF_X al_cc0b1799 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[45]));
  AL_DFF_X al_cc219e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a5e9c08d[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_930eb7ed[46]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_be310dbe (
    .a(1'b0),
    .o({al_50a889e9,open_n128}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d32d741c (
    .a(al_57dc9b0c[16]),
    .b(al_a5e9c08d[16]),
    .c(al_50a889e9),
    .o({al_45125ed0,al_d8106c92[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_14b2189d (
    .a(al_57dc9b0c[17]),
    .b(al_a5e9c08d[17]),
    .c(al_45125ed0),
    .o({al_256e1d30,al_d8106c92[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff04eb16 (
    .a(al_57dc9b0c[18]),
    .b(al_a5e9c08d[18]),
    .c(al_256e1d30),
    .o({al_6b8e1d26,al_d8106c92[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_810fbe40 (
    .a(al_57dc9b0c[19]),
    .b(al_a5e9c08d[19]),
    .c(al_6b8e1d26),
    .o({al_b57afe80,al_d8106c92[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ede5f176 (
    .a(al_57dc9b0c[20]),
    .b(al_a5e9c08d[20]),
    .c(al_b57afe80),
    .o({al_34a605a,al_d8106c92[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a82033e5 (
    .a(al_57dc9b0c[21]),
    .b(al_a5e9c08d[21]),
    .c(al_34a605a),
    .o({al_56bd060e,al_d8106c92[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_584f5d09 (
    .a(al_57dc9b0c[22]),
    .b(al_a5e9c08d[22]),
    .c(al_56bd060e),
    .o({al_c328a853,al_d8106c92[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_88fcb3bb (
    .a(al_57dc9b0c[23]),
    .b(al_a5e9c08d[23]),
    .c(al_c328a853),
    .o({al_4ffec454,al_d8106c92[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e98f2422 (
    .a(al_57dc9b0c[24]),
    .b(al_a5e9c08d[24]),
    .c(al_4ffec454),
    .o({al_d37de394,al_d8106c92[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_41b8ace3 (
    .a(al_57dc9b0c[25]),
    .b(al_a5e9c08d[25]),
    .c(al_d37de394),
    .o({al_1b2a14dc,al_d8106c92[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5ae00d90 (
    .a(al_57dc9b0c[26]),
    .b(al_a5e9c08d[26]),
    .c(al_1b2a14dc),
    .o({al_31a7b4b6,al_d8106c92[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ca6b00bd (
    .a(al_57dc9b0c[27]),
    .b(al_a5e9c08d[27]),
    .c(al_31a7b4b6),
    .o({al_d2a76de7,al_d8106c92[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b73a56c8 (
    .a(al_57dc9b0c[28]),
    .b(al_a5e9c08d[28]),
    .c(al_d2a76de7),
    .o({al_53f78588,al_d8106c92[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_277b5a62 (
    .a(al_57dc9b0c[29]),
    .b(al_a5e9c08d[29]),
    .c(al_53f78588),
    .o({al_89b70b3b,al_d8106c92[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_42f7b1c2 (
    .a(al_57dc9b0c[30]),
    .b(al_a5e9c08d[30]),
    .c(al_89b70b3b),
    .o({al_15cd8a93,al_d8106c92[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2a38efc7 (
    .a(al_57dc9b0c[31]),
    .b(al_a5e9c08d[31]),
    .c(al_15cd8a93),
    .o({al_eb481677,al_d8106c92[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3b44c2a4 (
    .a(al_57dc9b0c[32]),
    .b(al_a5e9c08d[32]),
    .c(al_eb481677),
    .o({al_1b3445fd,al_d8106c92[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dbe2453e (
    .a(al_57dc9b0c[33]),
    .b(al_a5e9c08d[33]),
    .c(al_1b3445fd),
    .o({al_1ab93794,al_d8106c92[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e8da2cd0 (
    .a(al_57dc9b0c[34]),
    .b(al_a5e9c08d[34]),
    .c(al_1ab93794),
    .o({al_c1f5ea1e,al_d8106c92[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_55c13538 (
    .a(al_57dc9b0c[35]),
    .b(al_a5e9c08d[35]),
    .c(al_c1f5ea1e),
    .o({al_57899523,al_d8106c92[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b67ffa21 (
    .a(al_57dc9b0c[36]),
    .b(al_a5e9c08d[36]),
    .c(al_57899523),
    .o({al_94297415,al_d8106c92[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d1e678c9 (
    .a(al_57dc9b0c[37]),
    .b(al_a5e9c08d[37]),
    .c(al_94297415),
    .o({al_1f080dc4,al_d8106c92[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_95bec237 (
    .a(al_57dc9b0c[38]),
    .b(al_a5e9c08d[38]),
    .c(al_1f080dc4),
    .o({al_de10dc85,al_d8106c92[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d5c95968 (
    .a(al_57dc9b0c[39]),
    .b(al_a5e9c08d[39]),
    .c(al_de10dc85),
    .o({al_b42d0d53,al_d8106c92[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ddab902 (
    .a(al_57dc9b0c[40]),
    .b(al_a5e9c08d[40]),
    .c(al_b42d0d53),
    .o({al_fd6c2091,al_d8106c92[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_415e46d6 (
    .a(al_57dc9b0c[41]),
    .b(al_a5e9c08d[41]),
    .c(al_fd6c2091),
    .o({al_c10da5dd,al_d8106c92[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3f8fb710 (
    .a(al_57dc9b0c[42]),
    .b(al_a5e9c08d[42]),
    .c(al_c10da5dd),
    .o({al_dd5f2a54,al_d8106c92[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f71fca3f (
    .a(al_57dc9b0c[43]),
    .b(al_a5e9c08d[43]),
    .c(al_dd5f2a54),
    .o({al_11eefeb5,al_d8106c92[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_134fd1f9 (
    .a(al_57dc9b0c[44]),
    .b(al_a5e9c08d[44]),
    .c(al_11eefeb5),
    .o({al_64eb948d,al_d8106c92[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_821b2144 (
    .a(al_57dc9b0c[45]),
    .b(al_a5e9c08d[45]),
    .c(al_64eb948d),
    .o({al_6ed7702d,al_d8106c92[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a4b3ec6 (
    .a(al_57dc9b0c[46]),
    .b(al_a5e9c08d[46]),
    .c(al_6ed7702d),
    .o({al_f68e810e,al_d8106c92[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a309e237 (
    .a(al_57dc9b0c[47]),
    .b(al_a5e9c08d[47]),
    .c(al_f68e810e),
    .o({al_430afd8b,al_d8106c92[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_99f2f050 (
    .a(1'b0),
    .b(1'b1),
    .c(al_430afd8b),
    .o({open_n129,al_f0ecaeb6}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_48654d0a (
    .a(al_57dc9b0c[16]),
    .b(al_d8106c92[0]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_42074f6b (
    .a(al_57dc9b0c[17]),
    .b(al_d8106c92[1]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9aaf0dc1 (
    .a(al_57dc9b0c[18]),
    .b(al_d8106c92[2]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8e71634d (
    .a(al_57dc9b0c[19]),
    .b(al_d8106c92[3]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6b7d1d91 (
    .a(al_57dc9b0c[20]),
    .b(al_d8106c92[4]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c4ca852d (
    .a(al_57dc9b0c[21]),
    .b(al_d8106c92[5]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4fbbad5a (
    .a(al_57dc9b0c[22]),
    .b(al_d8106c92[6]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9439a588 (
    .a(al_57dc9b0c[23]),
    .b(al_d8106c92[7]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_13239049 (
    .a(al_57dc9b0c[24]),
    .b(al_d8106c92[8]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1c4c4b16 (
    .a(al_57dc9b0c[25]),
    .b(al_d8106c92[9]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_84a0d2fc (
    .a(al_57dc9b0c[26]),
    .b(al_d8106c92[10]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f7fb8903 (
    .a(al_57dc9b0c[27]),
    .b(al_d8106c92[11]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_50f77443 (
    .a(al_57dc9b0c[28]),
    .b(al_d8106c92[12]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ae46e3e5 (
    .a(al_57dc9b0c[29]),
    .b(al_d8106c92[13]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ef45ea44 (
    .a(al_57dc9b0c[30]),
    .b(al_d8106c92[14]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_216990ac (
    .a(al_57dc9b0c[31]),
    .b(al_d8106c92[15]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cbf86a80 (
    .a(al_57dc9b0c[32]),
    .b(al_d8106c92[16]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_201e637f (
    .a(al_57dc9b0c[33]),
    .b(al_d8106c92[17]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_16928b24 (
    .a(al_57dc9b0c[34]),
    .b(al_d8106c92[18]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d52e7518 (
    .a(al_57dc9b0c[35]),
    .b(al_d8106c92[19]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b7dd4c02 (
    .a(al_57dc9b0c[36]),
    .b(al_d8106c92[20]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a87b7223 (
    .a(al_57dc9b0c[37]),
    .b(al_d8106c92[21]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_dfd792b3 (
    .a(al_57dc9b0c[38]),
    .b(al_d8106c92[22]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4aba126e (
    .a(al_57dc9b0c[39]),
    .b(al_d8106c92[23]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[39]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ca978822 (
    .a(al_57dc9b0c[40]),
    .b(al_d8106c92[24]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[40]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_35fd8d8 (
    .a(al_57dc9b0c[41]),
    .b(al_d8106c92[25]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[41]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9473b709 (
    .a(al_57dc9b0c[42]),
    .b(al_d8106c92[26]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[42]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ba94c099 (
    .a(al_57dc9b0c[43]),
    .b(al_d8106c92[27]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[43]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ac725169 (
    .a(al_57dc9b0c[44]),
    .b(al_d8106c92[28]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[44]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3ee62e3b (
    .a(al_57dc9b0c[45]),
    .b(al_d8106c92[29]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[45]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2d8d35b7 (
    .a(al_57dc9b0c[46]),
    .b(al_d8106c92[30]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[46]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_371330dc (
    .a(al_57dc9b0c[47]),
    .b(al_d8106c92[31]),
    .c(al_f0ecaeb6),
    .o(al_eb7d14b9[47]));
  AL_DFF_X al_3841317e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[0]));
  AL_DFF_X al_3a5017bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[9]));
  AL_DFF_X al_22bc7a0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[10]));
  AL_DFF_X al_3d8a9e16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[11]));
  AL_DFF_X al_81a57847 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[12]));
  AL_DFF_X al_ba2ccdd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[13]));
  AL_DFF_X al_830d689d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[14]));
  AL_DFF_X al_d18e6fbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[15]));
  AL_DFF_X al_cc948328 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[16]));
  AL_DFF_X al_b8068492 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[17]));
  AL_DFF_X al_3b38da80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[18]));
  AL_DFF_X al_e3c93dcf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[1]));
  AL_DFF_X al_a9ae3b5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[19]));
  AL_DFF_X al_fcd9c696 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[20]));
  AL_DFF_X al_a20b78a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[21]));
  AL_DFF_X al_8b043474 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[22]));
  AL_DFF_X al_1711d00e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[23]));
  AL_DFF_X al_d6eda739 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[24]));
  AL_DFF_X al_182d401 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[25]));
  AL_DFF_X al_e3f0c807 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[26]));
  AL_DFF_X al_3ef98cea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[27]));
  AL_DFF_X al_4696e9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[28]));
  AL_DFF_X al_2d9fa233 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[2]));
  AL_DFF_X al_f28d4341 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[29]));
  AL_DFF_X al_1c0e56f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[30]));
  AL_DFF_X al_e8321ef3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[31]));
  AL_DFF_X al_71e162be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[32]));
  AL_DFF_X al_4f729e7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[33]));
  AL_DFF_X al_f7fbceb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[34]));
  AL_DFF_X al_d9795af2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[35]));
  AL_DFF_X al_9b04d431 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[36]));
  AL_DFF_X al_cca9ebb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[37]));
  AL_DFF_X al_4e45a03a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[38]));
  AL_DFF_X al_c5f7cc67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[3]));
  AL_DFF_X al_29dea8db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[39]));
  AL_DFF_X al_d9e629ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[40]));
  AL_DFF_X al_6afdcbf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[41]));
  AL_DFF_X al_6dd696d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[42]));
  AL_DFF_X al_33847383 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[43]));
  AL_DFF_X al_50cc038e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[44]));
  AL_DFF_X al_c027db68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[45]));
  AL_DFF_X al_e4ed5b43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[46]));
  AL_DFF_X al_db825058 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_eb7d14b9[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[47]));
  AL_DFF_X al_cf65488d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[4]));
  AL_DFF_X al_8fd8c814 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[5]));
  AL_DFF_X al_d53e9d21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[6]));
  AL_DFF_X al_d72841e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[7]));
  AL_DFF_X al_e03e0796 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_57dc9b0c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_e7fdd367[8]));
  AL_DFF_X al_d4dc54a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f0ecaeb6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[0]));
  AL_DFF_X al_1fb097e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[9]));
  AL_DFF_X al_a3872f4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[10]));
  AL_DFF_X al_c6269498 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[11]));
  AL_DFF_X al_8fd7a822 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[12]));
  AL_DFF_X al_5fb31403 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[13]));
  AL_DFF_X al_f6748c30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[14]));
  AL_DFF_X al_71059bea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[15]));
  AL_DFF_X al_c71122d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[16]));
  AL_DFF_X al_17c252ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[17]));
  AL_DFF_X al_f78a85fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[18]));
  AL_DFF_X al_a3dc3707 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[1]));
  AL_DFF_X al_a10e26d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[19]));
  AL_DFF_X al_5d662ca0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[20]));
  AL_DFF_X al_6ecd9462 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[21]));
  AL_DFF_X al_1df1adf9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[22]));
  AL_DFF_X al_ab2560d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[23]));
  AL_DFF_X al_f17462bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[24]));
  AL_DFF_X al_909a60a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[25]));
  AL_DFF_X al_d5891080 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[26]));
  AL_DFF_X al_7868b64f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[27]));
  AL_DFF_X al_9ab3e9d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[28]));
  AL_DFF_X al_7ce40d66 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[2]));
  AL_DFF_X al_78fa98ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[29]));
  AL_DFF_X al_c7b38ef3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[30]));
  AL_DFF_X al_bac91f64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[31]));
  AL_DFF_X al_f80e262f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[3]));
  AL_DFF_X al_65618db5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[4]));
  AL_DFF_X al_6b94445d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[5]));
  AL_DFF_X al_5f183d8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[6]));
  AL_DFF_X al_fd400cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[7]));
  AL_DFF_X al_2aca26a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b40233aa[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_586198c7[8]));
  AL_DFF_X al_583c83d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2e2a074f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ad601da1[0]));
  AL_DFF_X al_a6fce482 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[14]));
  AL_DFF_X al_6704e0e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[15]));
  AL_DFF_X al_ce8f32ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[16]));
  AL_DFF_X al_fb22375 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[17]));
  AL_DFF_X al_a1803547 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[18]));
  AL_DFF_X al_6c2dca96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[19]));
  AL_DFF_X al_2318b073 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[20]));
  AL_DFF_X al_4e6e7e4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[21]));
  AL_DFF_X al_37991b0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[22]));
  AL_DFF_X al_c82fa9ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[23]));
  AL_DFF_X al_47e2a571 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[24]));
  AL_DFF_X al_28d7487e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[25]));
  AL_DFF_X al_52f0b5d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[26]));
  AL_DFF_X al_8d135949 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[27]));
  AL_DFF_X al_46d5b58b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[28]));
  AL_DFF_X al_a0cf4cfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[29]));
  AL_DFF_X al_5e01c96e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[30]));
  AL_DFF_X al_2d60263 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[31]));
  AL_DFF_X al_df56466c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[32]));
  AL_DFF_X al_294e1ed9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[33]));
  AL_DFF_X al_4dfe10e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[34]));
  AL_DFF_X al_90dab106 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[35]));
  AL_DFF_X al_95c22266 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[36]));
  AL_DFF_X al_3120a799 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[37]));
  AL_DFF_X al_300ddcb1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[38]));
  AL_DFF_X al_d10b4b54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[39]));
  AL_DFF_X al_5a0cb715 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[40]));
  AL_DFF_X al_cf9fd489 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[41]));
  AL_DFF_X al_2c94eb1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[42]));
  AL_DFF_X al_a6b4b66d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[43]));
  AL_DFF_X al_d14526f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[44]));
  AL_DFF_X al_8d2774c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_930eb7ed[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_400c3c08[45]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_a239d3a4 (
    .a(1'b0),
    .o({al_1376bcb0,open_n132}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b992ee2 (
    .a(al_e7fdd367[15]),
    .b(al_930eb7ed[15]),
    .c(al_1376bcb0),
    .o({al_4a06e815,al_ede1be73[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c31cb97e (
    .a(al_e7fdd367[16]),
    .b(al_930eb7ed[16]),
    .c(al_4a06e815),
    .o({al_58a18b68,al_ede1be73[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_df95de55 (
    .a(al_e7fdd367[17]),
    .b(al_930eb7ed[17]),
    .c(al_58a18b68),
    .o({al_4085a271,al_ede1be73[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2207a957 (
    .a(al_e7fdd367[18]),
    .b(al_930eb7ed[18]),
    .c(al_4085a271),
    .o({al_858f1c0c,al_ede1be73[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e104723d (
    .a(al_e7fdd367[19]),
    .b(al_930eb7ed[19]),
    .c(al_858f1c0c),
    .o({al_364abc0a,al_ede1be73[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_54f051be (
    .a(al_e7fdd367[20]),
    .b(al_930eb7ed[20]),
    .c(al_364abc0a),
    .o({al_9909f3ca,al_ede1be73[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2ea89ae2 (
    .a(al_e7fdd367[21]),
    .b(al_930eb7ed[21]),
    .c(al_9909f3ca),
    .o({al_bacdad1b,al_ede1be73[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_75463ff7 (
    .a(al_e7fdd367[22]),
    .b(al_930eb7ed[22]),
    .c(al_bacdad1b),
    .o({al_9bec1f33,al_ede1be73[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fec28a1d (
    .a(al_e7fdd367[23]),
    .b(al_930eb7ed[23]),
    .c(al_9bec1f33),
    .o({al_83f595b,al_ede1be73[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_16cbf829 (
    .a(al_e7fdd367[24]),
    .b(al_930eb7ed[24]),
    .c(al_83f595b),
    .o({al_91824dca,al_ede1be73[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a3ae4886 (
    .a(al_e7fdd367[25]),
    .b(al_930eb7ed[25]),
    .c(al_91824dca),
    .o({al_9ba07719,al_ede1be73[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e954911c (
    .a(al_e7fdd367[26]),
    .b(al_930eb7ed[26]),
    .c(al_9ba07719),
    .o({al_fc839793,al_ede1be73[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_160ad8ba (
    .a(al_e7fdd367[27]),
    .b(al_930eb7ed[27]),
    .c(al_fc839793),
    .o({al_739af9ca,al_ede1be73[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4ddc5cca (
    .a(al_e7fdd367[28]),
    .b(al_930eb7ed[28]),
    .c(al_739af9ca),
    .o({al_de14f218,al_ede1be73[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7aed9cc5 (
    .a(al_e7fdd367[29]),
    .b(al_930eb7ed[29]),
    .c(al_de14f218),
    .o({al_112db54d,al_ede1be73[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b232bafb (
    .a(al_e7fdd367[30]),
    .b(al_930eb7ed[30]),
    .c(al_112db54d),
    .o({al_f31a4cd8,al_ede1be73[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_99d0f9d1 (
    .a(al_e7fdd367[31]),
    .b(al_930eb7ed[31]),
    .c(al_f31a4cd8),
    .o({al_a77da9ed,al_ede1be73[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ee199cb7 (
    .a(al_e7fdd367[32]),
    .b(al_930eb7ed[32]),
    .c(al_a77da9ed),
    .o({al_9d63b53d,al_ede1be73[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_97f22f78 (
    .a(al_e7fdd367[33]),
    .b(al_930eb7ed[33]),
    .c(al_9d63b53d),
    .o({al_b187ff7c,al_ede1be73[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4a281389 (
    .a(al_e7fdd367[34]),
    .b(al_930eb7ed[34]),
    .c(al_b187ff7c),
    .o({al_a416feb9,al_ede1be73[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_25db82cd (
    .a(al_e7fdd367[35]),
    .b(al_930eb7ed[35]),
    .c(al_a416feb9),
    .o({al_3a2fee85,al_ede1be73[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4858fa5c (
    .a(al_e7fdd367[36]),
    .b(al_930eb7ed[36]),
    .c(al_3a2fee85),
    .o({al_af90c070,al_ede1be73[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3752267 (
    .a(al_e7fdd367[37]),
    .b(al_930eb7ed[37]),
    .c(al_af90c070),
    .o({al_a9f17098,al_ede1be73[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_28911eb7 (
    .a(al_e7fdd367[38]),
    .b(al_930eb7ed[38]),
    .c(al_a9f17098),
    .o({al_7b8d96e2,al_ede1be73[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dd71ef71 (
    .a(al_e7fdd367[39]),
    .b(al_930eb7ed[39]),
    .c(al_7b8d96e2),
    .o({al_a5b3371d,al_ede1be73[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_80e83d43 (
    .a(al_e7fdd367[40]),
    .b(al_930eb7ed[40]),
    .c(al_a5b3371d),
    .o({al_aa3a575d,al_ede1be73[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_922f4e6c (
    .a(al_e7fdd367[41]),
    .b(al_930eb7ed[41]),
    .c(al_aa3a575d),
    .o({al_354eea5a,al_ede1be73[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4c3f475d (
    .a(al_e7fdd367[42]),
    .b(al_930eb7ed[42]),
    .c(al_354eea5a),
    .o({al_94b0c7d1,al_ede1be73[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7ee9ae3e (
    .a(al_e7fdd367[43]),
    .b(al_930eb7ed[43]),
    .c(al_94b0c7d1),
    .o({al_cbca04a4,al_ede1be73[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b920650f (
    .a(al_e7fdd367[44]),
    .b(al_930eb7ed[44]),
    .c(al_cbca04a4),
    .o({al_9767aad8,al_ede1be73[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b37beab4 (
    .a(al_e7fdd367[45]),
    .b(al_930eb7ed[45]),
    .c(al_9767aad8),
    .o({al_1fe3c2d1,al_ede1be73[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_31488aa5 (
    .a(al_e7fdd367[46]),
    .b(al_930eb7ed[46]),
    .c(al_1fe3c2d1),
    .o({al_b233479,al_ede1be73[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_73c4d2bd (
    .a(al_e7fdd367[47]),
    .b(1'b0),
    .c(al_b233479),
    .o({al_71be4cd6,open_n133}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2fa8c8a1 (
    .a(1'b0),
    .b(1'b1),
    .c(al_71be4cd6),
    .o({open_n134,al_54a79559}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ee00f5a (
    .a(al_e7fdd367[15]),
    .b(al_ede1be73[0]),
    .c(al_54a79559),
    .o(al_f100da9b[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_787f4e8d (
    .a(al_e7fdd367[16]),
    .b(al_ede1be73[1]),
    .c(al_54a79559),
    .o(al_f100da9b[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a054920f (
    .a(al_e7fdd367[17]),
    .b(al_ede1be73[2]),
    .c(al_54a79559),
    .o(al_f100da9b[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1699698e (
    .a(al_e7fdd367[18]),
    .b(al_ede1be73[3]),
    .c(al_54a79559),
    .o(al_f100da9b[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b162044f (
    .a(al_e7fdd367[19]),
    .b(al_ede1be73[4]),
    .c(al_54a79559),
    .o(al_f100da9b[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9e1778d1 (
    .a(al_e7fdd367[20]),
    .b(al_ede1be73[5]),
    .c(al_54a79559),
    .o(al_f100da9b[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_eec7006c (
    .a(al_e7fdd367[21]),
    .b(al_ede1be73[6]),
    .c(al_54a79559),
    .o(al_f100da9b[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_747b45b0 (
    .a(al_e7fdd367[22]),
    .b(al_ede1be73[7]),
    .c(al_54a79559),
    .o(al_f100da9b[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_87438b1d (
    .a(al_e7fdd367[23]),
    .b(al_ede1be73[8]),
    .c(al_54a79559),
    .o(al_f100da9b[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_70d8f594 (
    .a(al_e7fdd367[24]),
    .b(al_ede1be73[9]),
    .c(al_54a79559),
    .o(al_f100da9b[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3ddbf56a (
    .a(al_e7fdd367[25]),
    .b(al_ede1be73[10]),
    .c(al_54a79559),
    .o(al_f100da9b[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b3595efa (
    .a(al_e7fdd367[26]),
    .b(al_ede1be73[11]),
    .c(al_54a79559),
    .o(al_f100da9b[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_90500fa5 (
    .a(al_e7fdd367[27]),
    .b(al_ede1be73[12]),
    .c(al_54a79559),
    .o(al_f100da9b[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a3bfc937 (
    .a(al_e7fdd367[28]),
    .b(al_ede1be73[13]),
    .c(al_54a79559),
    .o(al_f100da9b[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e836dc58 (
    .a(al_e7fdd367[29]),
    .b(al_ede1be73[14]),
    .c(al_54a79559),
    .o(al_f100da9b[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ce720c40 (
    .a(al_e7fdd367[30]),
    .b(al_ede1be73[15]),
    .c(al_54a79559),
    .o(al_f100da9b[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bba68974 (
    .a(al_e7fdd367[31]),
    .b(al_ede1be73[16]),
    .c(al_54a79559),
    .o(al_f100da9b[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d85460e1 (
    .a(al_e7fdd367[32]),
    .b(al_ede1be73[17]),
    .c(al_54a79559),
    .o(al_f100da9b[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_88cc63a6 (
    .a(al_e7fdd367[33]),
    .b(al_ede1be73[18]),
    .c(al_54a79559),
    .o(al_f100da9b[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_88e6e1d8 (
    .a(al_e7fdd367[34]),
    .b(al_ede1be73[19]),
    .c(al_54a79559),
    .o(al_f100da9b[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5dcfd5aa (
    .a(al_e7fdd367[35]),
    .b(al_ede1be73[20]),
    .c(al_54a79559),
    .o(al_f100da9b[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_37230d2a (
    .a(al_e7fdd367[36]),
    .b(al_ede1be73[21]),
    .c(al_54a79559),
    .o(al_f100da9b[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_be9be112 (
    .a(al_e7fdd367[37]),
    .b(al_ede1be73[22]),
    .c(al_54a79559),
    .o(al_f100da9b[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_41b60aa7 (
    .a(al_e7fdd367[38]),
    .b(al_ede1be73[23]),
    .c(al_54a79559),
    .o(al_f100da9b[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_431227bb (
    .a(al_e7fdd367[39]),
    .b(al_ede1be73[24]),
    .c(al_54a79559),
    .o(al_f100da9b[39]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_389916c6 (
    .a(al_e7fdd367[40]),
    .b(al_ede1be73[25]),
    .c(al_54a79559),
    .o(al_f100da9b[40]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b4cbcee7 (
    .a(al_e7fdd367[41]),
    .b(al_ede1be73[26]),
    .c(al_54a79559),
    .o(al_f100da9b[41]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2c089c6 (
    .a(al_e7fdd367[42]),
    .b(al_ede1be73[27]),
    .c(al_54a79559),
    .o(al_f100da9b[42]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a5e30c4f (
    .a(al_e7fdd367[43]),
    .b(al_ede1be73[28]),
    .c(al_54a79559),
    .o(al_f100da9b[43]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_50a3607a (
    .a(al_e7fdd367[44]),
    .b(al_ede1be73[29]),
    .c(al_54a79559),
    .o(al_f100da9b[44]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c4199fcb (
    .a(al_e7fdd367[45]),
    .b(al_ede1be73[30]),
    .c(al_54a79559),
    .o(al_f100da9b[45]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5f52ba78 (
    .a(al_e7fdd367[46]),
    .b(al_ede1be73[31]),
    .c(al_54a79559),
    .o(al_f100da9b[46]));
  AL_DFF_X al_84722c1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[0]));
  AL_DFF_X al_ef1801f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[9]));
  AL_DFF_X al_bdb21074 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[10]));
  AL_DFF_X al_c012de4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[11]));
  AL_DFF_X al_374c89a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[12]));
  AL_DFF_X al_6b446070 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[13]));
  AL_DFF_X al_a97079a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[14]));
  AL_DFF_X al_1e6a2d01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[15]));
  AL_DFF_X al_298b323f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[16]));
  AL_DFF_X al_c29ea134 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[17]));
  AL_DFF_X al_b1a32edf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[18]));
  AL_DFF_X al_71483aba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[1]));
  AL_DFF_X al_a19331ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[19]));
  AL_DFF_X al_479bef7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[20]));
  AL_DFF_X al_941e5ae3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[21]));
  AL_DFF_X al_41f5ec1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[22]));
  AL_DFF_X al_16fbda (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[23]));
  AL_DFF_X al_f914b0f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[24]));
  AL_DFF_X al_9df8a449 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[25]));
  AL_DFF_X al_2093bccc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[26]));
  AL_DFF_X al_842a2e26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[27]));
  AL_DFF_X al_8a90562c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[28]));
  AL_DFF_X al_8e1dc2a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[2]));
  AL_DFF_X al_2fdb95e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[29]));
  AL_DFF_X al_1fb3ed0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[30]));
  AL_DFF_X al_b33554e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[31]));
  AL_DFF_X al_d2603c07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[32]));
  AL_DFF_X al_8d5a165a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[33]));
  AL_DFF_X al_ba0f3baa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[34]));
  AL_DFF_X al_5f2d088 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[35]));
  AL_DFF_X al_84300af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[36]));
  AL_DFF_X al_b8d7e51d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[37]));
  AL_DFF_X al_566ac786 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[38]));
  AL_DFF_X al_465ee902 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[3]));
  AL_DFF_X al_88b7b46e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[39]));
  AL_DFF_X al_413fd5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[40]));
  AL_DFF_X al_49193e1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[41]));
  AL_DFF_X al_fadb6797 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[42]));
  AL_DFF_X al_21939527 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[43]));
  AL_DFF_X al_87418710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[44]));
  AL_DFF_X al_b3f6df7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[45]));
  AL_DFF_X al_be609446 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f100da9b[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[46]));
  AL_DFF_X al_83aef2ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[4]));
  AL_DFF_X al_97f76716 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[5]));
  AL_DFF_X al_eea9357 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[6]));
  AL_DFF_X al_c7b9b3f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[7]));
  AL_DFF_X al_316cfdd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e7fdd367[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5675a322[8]));
  AL_DFF_X al_e44aa87f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_54a79559),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[0]));
  AL_DFF_X al_18f8c396 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[9]));
  AL_DFF_X al_d479ff4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[10]));
  AL_DFF_X al_38136589 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[11]));
  AL_DFF_X al_c37df49b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[12]));
  AL_DFF_X al_89e5a599 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[13]));
  AL_DFF_X al_8ff8fb72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[14]));
  AL_DFF_X al_9e170378 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[15]));
  AL_DFF_X al_97c75b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[16]));
  AL_DFF_X al_f9dd3c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[17]));
  AL_DFF_X al_9c13ad60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[18]));
  AL_DFF_X al_e7a631d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[1]));
  AL_DFF_X al_ae205687 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[19]));
  AL_DFF_X al_73107ead (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[20]));
  AL_DFF_X al_8238c2da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[21]));
  AL_DFF_X al_46bcc6b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[22]));
  AL_DFF_X al_d11b642e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[23]));
  AL_DFF_X al_641e06ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[24]));
  AL_DFF_X al_fbac7fc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[25]));
  AL_DFF_X al_83dd9bd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[26]));
  AL_DFF_X al_d12a6508 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[27]));
  AL_DFF_X al_ce15a3c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[28]));
  AL_DFF_X al_103d9b82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[2]));
  AL_DFF_X al_9b210777 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[29]));
  AL_DFF_X al_1f903cb3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[30]));
  AL_DFF_X al_31a2467b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[31]));
  AL_DFF_X al_cf2f7566 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[32]));
  AL_DFF_X al_d1677d83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[3]));
  AL_DFF_X al_4411b2a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[4]));
  AL_DFF_X al_f34b89fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[5]));
  AL_DFF_X al_1357e6dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[6]));
  AL_DFF_X al_8414ffda (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[7]));
  AL_DFF_X al_8cd0a95f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_586198c7[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3a0a3044[8]));
  AL_DFF_X al_f79f51db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ad601da1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ff0af5c2[0]));
  AL_DFF_X al_c9a1c844 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[13]));
  AL_DFF_X al_16397e6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[14]));
  AL_DFF_X al_f017a78c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[15]));
  AL_DFF_X al_5fc19ff3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[16]));
  AL_DFF_X al_225ffe6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[17]));
  AL_DFF_X al_f5957a9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[18]));
  AL_DFF_X al_4f7f04a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[19]));
  AL_DFF_X al_53423d56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[20]));
  AL_DFF_X al_cf8a1668 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[21]));
  AL_DFF_X al_641c66df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[22]));
  AL_DFF_X al_67e9ca36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[23]));
  AL_DFF_X al_a191918f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[24]));
  AL_DFF_X al_bb1193ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[25]));
  AL_DFF_X al_de454188 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[26]));
  AL_DFF_X al_5bfd2703 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[27]));
  AL_DFF_X al_b84bdf4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[28]));
  AL_DFF_X al_8c2df796 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[29]));
  AL_DFF_X al_10fd89d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[30]));
  AL_DFF_X al_58d5c88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[31]));
  AL_DFF_X al_6cd81b72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[32]));
  AL_DFF_X al_a4919633 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[33]));
  AL_DFF_X al_a27600ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[34]));
  AL_DFF_X al_ab816685 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[35]));
  AL_DFF_X al_99974655 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[36]));
  AL_DFF_X al_347e41b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[37]));
  AL_DFF_X al_8780814e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[38]));
  AL_DFF_X al_410a29a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[39]));
  AL_DFF_X al_c2d5dcb4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[40]));
  AL_DFF_X al_4268fba9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[41]));
  AL_DFF_X al_7b5b36aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[42]));
  AL_DFF_X al_c8ba2ce1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[43]));
  AL_DFF_X al_b8ec4bed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_400c3c08[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_304b2866[44]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_289d9316 (
    .a(1'b0),
    .o({al_c4782520,open_n137}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c9d4554a (
    .a(al_5675a322[14]),
    .b(al_400c3c08[14]),
    .c(al_c4782520),
    .o({al_b1f716e3,al_2232b9e8[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b7744df3 (
    .a(al_5675a322[15]),
    .b(al_400c3c08[15]),
    .c(al_b1f716e3),
    .o({al_a59de26c,al_2232b9e8[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f8d6524a (
    .a(al_5675a322[16]),
    .b(al_400c3c08[16]),
    .c(al_a59de26c),
    .o({al_561ce4c4,al_2232b9e8[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_97332442 (
    .a(al_5675a322[17]),
    .b(al_400c3c08[17]),
    .c(al_561ce4c4),
    .o({al_2451e527,al_2232b9e8[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_829251c9 (
    .a(al_5675a322[18]),
    .b(al_400c3c08[18]),
    .c(al_2451e527),
    .o({al_2bed1d6f,al_2232b9e8[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9d7b018a (
    .a(al_5675a322[19]),
    .b(al_400c3c08[19]),
    .c(al_2bed1d6f),
    .o({al_a9898f67,al_2232b9e8[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_50834aaf (
    .a(al_5675a322[20]),
    .b(al_400c3c08[20]),
    .c(al_a9898f67),
    .o({al_7999a920,al_2232b9e8[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b35c65b6 (
    .a(al_5675a322[21]),
    .b(al_400c3c08[21]),
    .c(al_7999a920),
    .o({al_dcd3196f,al_2232b9e8[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e912a8a4 (
    .a(al_5675a322[22]),
    .b(al_400c3c08[22]),
    .c(al_dcd3196f),
    .o({al_9d1db55,al_2232b9e8[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_163687c8 (
    .a(al_5675a322[23]),
    .b(al_400c3c08[23]),
    .c(al_9d1db55),
    .o({al_9240c8a4,al_2232b9e8[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e562e65f (
    .a(al_5675a322[24]),
    .b(al_400c3c08[24]),
    .c(al_9240c8a4),
    .o({al_f5953bb1,al_2232b9e8[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9cbc3de8 (
    .a(al_5675a322[25]),
    .b(al_400c3c08[25]),
    .c(al_f5953bb1),
    .o({al_ff96e0f,al_2232b9e8[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40945769 (
    .a(al_5675a322[26]),
    .b(al_400c3c08[26]),
    .c(al_ff96e0f),
    .o({al_fdc157ff,al_2232b9e8[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_26251102 (
    .a(al_5675a322[27]),
    .b(al_400c3c08[27]),
    .c(al_fdc157ff),
    .o({al_fa3f4f58,al_2232b9e8[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6f354661 (
    .a(al_5675a322[28]),
    .b(al_400c3c08[28]),
    .c(al_fa3f4f58),
    .o({al_f0643c82,al_2232b9e8[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2ab19757 (
    .a(al_5675a322[29]),
    .b(al_400c3c08[29]),
    .c(al_f0643c82),
    .o({al_1106f695,al_2232b9e8[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_504577a6 (
    .a(al_5675a322[30]),
    .b(al_400c3c08[30]),
    .c(al_1106f695),
    .o({al_474d64a7,al_2232b9e8[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1fa0565f (
    .a(al_5675a322[31]),
    .b(al_400c3c08[31]),
    .c(al_474d64a7),
    .o({al_d079fcc4,al_2232b9e8[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1d988baf (
    .a(al_5675a322[32]),
    .b(al_400c3c08[32]),
    .c(al_d079fcc4),
    .o({al_8af08334,al_2232b9e8[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_59e6b8ba (
    .a(al_5675a322[33]),
    .b(al_400c3c08[33]),
    .c(al_8af08334),
    .o({al_d3786c88,al_2232b9e8[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4b42c71b (
    .a(al_5675a322[34]),
    .b(al_400c3c08[34]),
    .c(al_d3786c88),
    .o({al_1c2d1a70,al_2232b9e8[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_82754b5b (
    .a(al_5675a322[35]),
    .b(al_400c3c08[35]),
    .c(al_1c2d1a70),
    .o({al_47dadb08,al_2232b9e8[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b550afa4 (
    .a(al_5675a322[36]),
    .b(al_400c3c08[36]),
    .c(al_47dadb08),
    .o({al_4145de8a,al_2232b9e8[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a8c2fd16 (
    .a(al_5675a322[37]),
    .b(al_400c3c08[37]),
    .c(al_4145de8a),
    .o({al_1dddd2e5,al_2232b9e8[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bf792b58 (
    .a(al_5675a322[38]),
    .b(al_400c3c08[38]),
    .c(al_1dddd2e5),
    .o({al_90ad6b5d,al_2232b9e8[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_70d52565 (
    .a(al_5675a322[39]),
    .b(al_400c3c08[39]),
    .c(al_90ad6b5d),
    .o({al_f4e9ff5b,al_2232b9e8[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_14dc5efc (
    .a(al_5675a322[40]),
    .b(al_400c3c08[40]),
    .c(al_f4e9ff5b),
    .o({al_615d34bc,al_2232b9e8[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_84a3a78 (
    .a(al_5675a322[41]),
    .b(al_400c3c08[41]),
    .c(al_615d34bc),
    .o({al_7b56c629,al_2232b9e8[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cd43dde (
    .a(al_5675a322[42]),
    .b(al_400c3c08[42]),
    .c(al_7b56c629),
    .o({al_90865e32,al_2232b9e8[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a5f643b3 (
    .a(al_5675a322[43]),
    .b(al_400c3c08[43]),
    .c(al_90865e32),
    .o({al_5bc29d76,al_2232b9e8[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1c5128d6 (
    .a(al_5675a322[44]),
    .b(al_400c3c08[44]),
    .c(al_5bc29d76),
    .o({al_b89115b,al_2232b9e8[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c7397a60 (
    .a(al_5675a322[45]),
    .b(al_400c3c08[45]),
    .c(al_b89115b),
    .o({al_1bed3aa5,al_2232b9e8[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3c6ae6b0 (
    .a(al_5675a322[46]),
    .b(1'b0),
    .c(al_1bed3aa5),
    .o({al_ee91a42b,open_n138}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b76d295b (
    .a(1'b0),
    .b(1'b1),
    .c(al_ee91a42b),
    .o({open_n139,al_d9039a1f}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_17e70baf (
    .a(al_5675a322[14]),
    .b(al_2232b9e8[0]),
    .c(al_d9039a1f),
    .o(al_dacf1710[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ea5767db (
    .a(al_5675a322[15]),
    .b(al_2232b9e8[1]),
    .c(al_d9039a1f),
    .o(al_dacf1710[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_98a42982 (
    .a(al_5675a322[16]),
    .b(al_2232b9e8[2]),
    .c(al_d9039a1f),
    .o(al_dacf1710[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7557e1cc (
    .a(al_5675a322[17]),
    .b(al_2232b9e8[3]),
    .c(al_d9039a1f),
    .o(al_dacf1710[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2fe449e1 (
    .a(al_5675a322[18]),
    .b(al_2232b9e8[4]),
    .c(al_d9039a1f),
    .o(al_dacf1710[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_51f38d0c (
    .a(al_5675a322[19]),
    .b(al_2232b9e8[5]),
    .c(al_d9039a1f),
    .o(al_dacf1710[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_32e8d4b4 (
    .a(al_5675a322[20]),
    .b(al_2232b9e8[6]),
    .c(al_d9039a1f),
    .o(al_dacf1710[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_125ee0df (
    .a(al_5675a322[21]),
    .b(al_2232b9e8[7]),
    .c(al_d9039a1f),
    .o(al_dacf1710[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c61f2457 (
    .a(al_5675a322[22]),
    .b(al_2232b9e8[8]),
    .c(al_d9039a1f),
    .o(al_dacf1710[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4fd6094e (
    .a(al_5675a322[23]),
    .b(al_2232b9e8[9]),
    .c(al_d9039a1f),
    .o(al_dacf1710[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_61dae153 (
    .a(al_5675a322[24]),
    .b(al_2232b9e8[10]),
    .c(al_d9039a1f),
    .o(al_dacf1710[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_52e845aa (
    .a(al_5675a322[25]),
    .b(al_2232b9e8[11]),
    .c(al_d9039a1f),
    .o(al_dacf1710[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7ebeb00c (
    .a(al_5675a322[26]),
    .b(al_2232b9e8[12]),
    .c(al_d9039a1f),
    .o(al_dacf1710[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f088bed (
    .a(al_5675a322[27]),
    .b(al_2232b9e8[13]),
    .c(al_d9039a1f),
    .o(al_dacf1710[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1b70cb0f (
    .a(al_5675a322[28]),
    .b(al_2232b9e8[14]),
    .c(al_d9039a1f),
    .o(al_dacf1710[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ae687152 (
    .a(al_5675a322[29]),
    .b(al_2232b9e8[15]),
    .c(al_d9039a1f),
    .o(al_dacf1710[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fcec6549 (
    .a(al_5675a322[30]),
    .b(al_2232b9e8[16]),
    .c(al_d9039a1f),
    .o(al_dacf1710[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_33402414 (
    .a(al_5675a322[31]),
    .b(al_2232b9e8[17]),
    .c(al_d9039a1f),
    .o(al_dacf1710[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a9149aab (
    .a(al_5675a322[32]),
    .b(al_2232b9e8[18]),
    .c(al_d9039a1f),
    .o(al_dacf1710[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_743454da (
    .a(al_5675a322[33]),
    .b(al_2232b9e8[19]),
    .c(al_d9039a1f),
    .o(al_dacf1710[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8ea4d5bd (
    .a(al_5675a322[34]),
    .b(al_2232b9e8[20]),
    .c(al_d9039a1f),
    .o(al_dacf1710[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_43107c3d (
    .a(al_5675a322[35]),
    .b(al_2232b9e8[21]),
    .c(al_d9039a1f),
    .o(al_dacf1710[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b67d97dc (
    .a(al_5675a322[36]),
    .b(al_2232b9e8[22]),
    .c(al_d9039a1f),
    .o(al_dacf1710[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_efac167e (
    .a(al_5675a322[37]),
    .b(al_2232b9e8[23]),
    .c(al_d9039a1f),
    .o(al_dacf1710[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4bc8bb58 (
    .a(al_5675a322[38]),
    .b(al_2232b9e8[24]),
    .c(al_d9039a1f),
    .o(al_dacf1710[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9ad67346 (
    .a(al_5675a322[39]),
    .b(al_2232b9e8[25]),
    .c(al_d9039a1f),
    .o(al_dacf1710[39]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8e0bb556 (
    .a(al_5675a322[40]),
    .b(al_2232b9e8[26]),
    .c(al_d9039a1f),
    .o(al_dacf1710[40]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6c5e7e05 (
    .a(al_5675a322[41]),
    .b(al_2232b9e8[27]),
    .c(al_d9039a1f),
    .o(al_dacf1710[41]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_98155397 (
    .a(al_5675a322[42]),
    .b(al_2232b9e8[28]),
    .c(al_d9039a1f),
    .o(al_dacf1710[42]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7b6abcbb (
    .a(al_5675a322[43]),
    .b(al_2232b9e8[29]),
    .c(al_d9039a1f),
    .o(al_dacf1710[43]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_732b9be9 (
    .a(al_5675a322[44]),
    .b(al_2232b9e8[30]),
    .c(al_d9039a1f),
    .o(al_dacf1710[44]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_821bf45d (
    .a(al_5675a322[45]),
    .b(al_2232b9e8[31]),
    .c(al_d9039a1f),
    .o(al_dacf1710[45]));
  AL_DFF_X al_c8342c44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[0]));
  AL_DFF_X al_3b768ec2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[9]));
  AL_DFF_X al_ff3e335c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[10]));
  AL_DFF_X al_4063a59e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[11]));
  AL_DFF_X al_a12b6262 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[12]));
  AL_DFF_X al_562799da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[13]));
  AL_DFF_X al_1003a87a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[14]));
  AL_DFF_X al_ccf7c729 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[15]));
  AL_DFF_X al_cc131c14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[16]));
  AL_DFF_X al_bc18762c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[17]));
  AL_DFF_X al_2e5d32da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[18]));
  AL_DFF_X al_a47186ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[1]));
  AL_DFF_X al_1eab4aaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[19]));
  AL_DFF_X al_72859a52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[20]));
  AL_DFF_X al_13183806 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[21]));
  AL_DFF_X al_a8e099af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[22]));
  AL_DFF_X al_feab60b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[23]));
  AL_DFF_X al_dbdb465a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[24]));
  AL_DFF_X al_5c862336 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[25]));
  AL_DFF_X al_e5e84e34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[26]));
  AL_DFF_X al_784edc1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[27]));
  AL_DFF_X al_d211e782 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[28]));
  AL_DFF_X al_26655355 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[2]));
  AL_DFF_X al_b0a19bd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[29]));
  AL_DFF_X al_8660ca33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[30]));
  AL_DFF_X al_f5f6327a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[31]));
  AL_DFF_X al_4fa7d8df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[32]));
  AL_DFF_X al_392b1efa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[33]));
  AL_DFF_X al_34b61d4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[34]));
  AL_DFF_X al_2f7cbdfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[35]));
  AL_DFF_X al_5c51c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[36]));
  AL_DFF_X al_dec0126b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[37]));
  AL_DFF_X al_68d69e92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[38]));
  AL_DFF_X al_41b84fd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[3]));
  AL_DFF_X al_3abea39b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[39]));
  AL_DFF_X al_8afdffa5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[40]));
  AL_DFF_X al_2242bfac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[41]));
  AL_DFF_X al_48fc9890 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[42]));
  AL_DFF_X al_e0f74106 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[43]));
  AL_DFF_X al_17b65e5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[44]));
  AL_DFF_X al_433981ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dacf1710[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[45]));
  AL_DFF_X al_ff65032e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[4]));
  AL_DFF_X al_c6667dcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[5]));
  AL_DFF_X al_5b327aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[6]));
  AL_DFF_X al_d8133f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[7]));
  AL_DFF_X al_2cf505a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5675a322[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c7be2582[8]));
  AL_DFF_X al_222853c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9039a1f),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[0]));
  AL_DFF_X al_29e20947 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[9]));
  AL_DFF_X al_e9a586fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[10]));
  AL_DFF_X al_4171a53e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[11]));
  AL_DFF_X al_340ffc55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[12]));
  AL_DFF_X al_a16d2960 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[13]));
  AL_DFF_X al_d9c1f5c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[14]));
  AL_DFF_X al_81d6020f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[15]));
  AL_DFF_X al_9f2252eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[16]));
  AL_DFF_X al_5398c839 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[17]));
  AL_DFF_X al_ec64cd97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[18]));
  AL_DFF_X al_37ba6fdf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[1]));
  AL_DFF_X al_764241ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[19]));
  AL_DFF_X al_6d3f756f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[20]));
  AL_DFF_X al_3a2aae8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[21]));
  AL_DFF_X al_c94c2bdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[22]));
  AL_DFF_X al_1f44d37a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[23]));
  AL_DFF_X al_9e76919 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[24]));
  AL_DFF_X al_f5760323 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[25]));
  AL_DFF_X al_4559d368 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[26]));
  AL_DFF_X al_7b57cb1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[27]));
  AL_DFF_X al_22c2895b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[28]));
  AL_DFF_X al_d7d474c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[2]));
  AL_DFF_X al_5ff25236 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[29]));
  AL_DFF_X al_ac7f7d16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[30]));
  AL_DFF_X al_6dc46472 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[31]));
  AL_DFF_X al_f5c02724 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[32]));
  AL_DFF_X al_a5073be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[33]));
  AL_DFF_X al_754bd3a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[3]));
  AL_DFF_X al_ff7b2a84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[4]));
  AL_DFF_X al_3ffc0e82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[5]));
  AL_DFF_X al_edbd467b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[6]));
  AL_DFF_X al_6fe741ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[7]));
  AL_DFF_X al_8a3ad9fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3a0a3044[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_64e3fb17[8]));
  AL_DFF_X al_a623f572 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ff0af5c2[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_65c09044[0]));
  AL_DFF_X al_9168e28d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[12]));
  AL_DFF_X al_599651f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[13]));
  AL_DFF_X al_58aff662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[14]));
  AL_DFF_X al_eef52afb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[15]));
  AL_DFF_X al_1ccba987 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[16]));
  AL_DFF_X al_b78f42fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[17]));
  AL_DFF_X al_a320bd6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[18]));
  AL_DFF_X al_82ee14cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[19]));
  AL_DFF_X al_15a5c75e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[20]));
  AL_DFF_X al_34930d9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[21]));
  AL_DFF_X al_13670aca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[22]));
  AL_DFF_X al_8d6dc775 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[23]));
  AL_DFF_X al_8a019b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[24]));
  AL_DFF_X al_227ce989 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[25]));
  AL_DFF_X al_424888de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[26]));
  AL_DFF_X al_9567cf16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[27]));
  AL_DFF_X al_79e8091e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[28]));
  AL_DFF_X al_7040be7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[29]));
  AL_DFF_X al_47473e39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[30]));
  AL_DFF_X al_dd217966 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[31]));
  AL_DFF_X al_90b6633d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[32]));
  AL_DFF_X al_67e9b7da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[33]));
  AL_DFF_X al_73c578ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[34]));
  AL_DFF_X al_f75959f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[35]));
  AL_DFF_X al_c3b898fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[36]));
  AL_DFF_X al_3bf81386 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[37]));
  AL_DFF_X al_6f79341f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[38]));
  AL_DFF_X al_9b0c4091 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[39]));
  AL_DFF_X al_c908002c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[40]));
  AL_DFF_X al_a441a8cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[41]));
  AL_DFF_X al_5ade803 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[42]));
  AL_DFF_X al_9a21955c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_304b2866[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bac230e2[43]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_51b0a9ce (
    .a(1'b0),
    .o({al_5dced79d,open_n142}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_59b69438 (
    .a(al_c7be2582[13]),
    .b(al_304b2866[13]),
    .c(al_5dced79d),
    .o({al_c2c29ff3,al_fab6b65e[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_11ce12ad (
    .a(al_c7be2582[14]),
    .b(al_304b2866[14]),
    .c(al_c2c29ff3),
    .o({al_bb679170,al_fab6b65e[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e9001853 (
    .a(al_c7be2582[15]),
    .b(al_304b2866[15]),
    .c(al_bb679170),
    .o({al_e9214bad,al_fab6b65e[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_62a22ab0 (
    .a(al_c7be2582[16]),
    .b(al_304b2866[16]),
    .c(al_e9214bad),
    .o({al_a13e1232,al_fab6b65e[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5f77a2a7 (
    .a(al_c7be2582[17]),
    .b(al_304b2866[17]),
    .c(al_a13e1232),
    .o({al_e9639971,al_fab6b65e[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d61117ad (
    .a(al_c7be2582[18]),
    .b(al_304b2866[18]),
    .c(al_e9639971),
    .o({al_15e685d4,al_fab6b65e[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40dad8a2 (
    .a(al_c7be2582[19]),
    .b(al_304b2866[19]),
    .c(al_15e685d4),
    .o({al_d09dedfa,al_fab6b65e[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_928373a3 (
    .a(al_c7be2582[20]),
    .b(al_304b2866[20]),
    .c(al_d09dedfa),
    .o({al_d38c342e,al_fab6b65e[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4451110d (
    .a(al_c7be2582[21]),
    .b(al_304b2866[21]),
    .c(al_d38c342e),
    .o({al_718df034,al_fab6b65e[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d44ae6dd (
    .a(al_c7be2582[22]),
    .b(al_304b2866[22]),
    .c(al_718df034),
    .o({al_97f6d29,al_fab6b65e[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d4cd8f52 (
    .a(al_c7be2582[23]),
    .b(al_304b2866[23]),
    .c(al_97f6d29),
    .o({al_d87faa07,al_fab6b65e[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b76eef6b (
    .a(al_c7be2582[24]),
    .b(al_304b2866[24]),
    .c(al_d87faa07),
    .o({al_f45a16f4,al_fab6b65e[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_acd48e99 (
    .a(al_c7be2582[25]),
    .b(al_304b2866[25]),
    .c(al_f45a16f4),
    .o({al_23c32ed1,al_fab6b65e[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4d3123e6 (
    .a(al_c7be2582[26]),
    .b(al_304b2866[26]),
    .c(al_23c32ed1),
    .o({al_5c729632,al_fab6b65e[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b13eb446 (
    .a(al_c7be2582[27]),
    .b(al_304b2866[27]),
    .c(al_5c729632),
    .o({al_117d184b,al_fab6b65e[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7f0113ea (
    .a(al_c7be2582[28]),
    .b(al_304b2866[28]),
    .c(al_117d184b),
    .o({al_cd65094,al_fab6b65e[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f7887586 (
    .a(al_c7be2582[29]),
    .b(al_304b2866[29]),
    .c(al_cd65094),
    .o({al_cdc4fc2e,al_fab6b65e[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_83b4f2aa (
    .a(al_c7be2582[30]),
    .b(al_304b2866[30]),
    .c(al_cdc4fc2e),
    .o({al_88c69413,al_fab6b65e[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17061929 (
    .a(al_c7be2582[31]),
    .b(al_304b2866[31]),
    .c(al_88c69413),
    .o({al_624a5f2d,al_fab6b65e[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c0178d48 (
    .a(al_c7be2582[32]),
    .b(al_304b2866[32]),
    .c(al_624a5f2d),
    .o({al_d71b24d6,al_fab6b65e[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3fb7096b (
    .a(al_c7be2582[33]),
    .b(al_304b2866[33]),
    .c(al_d71b24d6),
    .o({al_a1d5dec3,al_fab6b65e[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_497b0f3a (
    .a(al_c7be2582[34]),
    .b(al_304b2866[34]),
    .c(al_a1d5dec3),
    .o({al_12dadb42,al_fab6b65e[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ac0f6ddd (
    .a(al_c7be2582[35]),
    .b(al_304b2866[35]),
    .c(al_12dadb42),
    .o({al_bc1185ef,al_fab6b65e[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc0f8fa2 (
    .a(al_c7be2582[36]),
    .b(al_304b2866[36]),
    .c(al_bc1185ef),
    .o({al_d5531fd2,al_fab6b65e[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a7da32de (
    .a(al_c7be2582[37]),
    .b(al_304b2866[37]),
    .c(al_d5531fd2),
    .o({al_b07fbb26,al_fab6b65e[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3e1b6ed0 (
    .a(al_c7be2582[38]),
    .b(al_304b2866[38]),
    .c(al_b07fbb26),
    .o({al_8a3c5223,al_fab6b65e[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_16f97b3d (
    .a(al_c7be2582[39]),
    .b(al_304b2866[39]),
    .c(al_8a3c5223),
    .o({al_4dd1780b,al_fab6b65e[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1701c4b0 (
    .a(al_c7be2582[40]),
    .b(al_304b2866[40]),
    .c(al_4dd1780b),
    .o({al_a06e1c18,al_fab6b65e[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_57b07e3e (
    .a(al_c7be2582[41]),
    .b(al_304b2866[41]),
    .c(al_a06e1c18),
    .o({al_50022df0,al_fab6b65e[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d1712071 (
    .a(al_c7be2582[42]),
    .b(al_304b2866[42]),
    .c(al_50022df0),
    .o({al_58ce9b0f,al_fab6b65e[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ad68580b (
    .a(al_c7be2582[43]),
    .b(al_304b2866[43]),
    .c(al_58ce9b0f),
    .o({al_542e503f,al_fab6b65e[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3c0aa229 (
    .a(al_c7be2582[44]),
    .b(al_304b2866[44]),
    .c(al_542e503f),
    .o({al_55bbc798,al_fab6b65e[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2bb3dd01 (
    .a(al_c7be2582[45]),
    .b(1'b0),
    .c(al_55bbc798),
    .o({al_aa5ae88a,open_n143}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc0dfd0f (
    .a(1'b0),
    .b(1'b1),
    .c(al_aa5ae88a),
    .o({open_n144,al_5b4dd00b}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_de302e73 (
    .a(al_c7be2582[13]),
    .b(al_fab6b65e[0]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e46899d5 (
    .a(al_c7be2582[14]),
    .b(al_fab6b65e[1]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6f03137a (
    .a(al_c7be2582[15]),
    .b(al_fab6b65e[2]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d2a486fa (
    .a(al_c7be2582[16]),
    .b(al_fab6b65e[3]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fc165eed (
    .a(al_c7be2582[17]),
    .b(al_fab6b65e[4]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8c2588ed (
    .a(al_c7be2582[18]),
    .b(al_fab6b65e[5]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6a28f135 (
    .a(al_c7be2582[19]),
    .b(al_fab6b65e[6]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5ca4f75d (
    .a(al_c7be2582[20]),
    .b(al_fab6b65e[7]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f1a9da2d (
    .a(al_c7be2582[21]),
    .b(al_fab6b65e[8]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bace43c (
    .a(al_c7be2582[22]),
    .b(al_fab6b65e[9]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bfec82ac (
    .a(al_c7be2582[23]),
    .b(al_fab6b65e[10]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a39f7dae (
    .a(al_c7be2582[24]),
    .b(al_fab6b65e[11]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_399a7d5d (
    .a(al_c7be2582[25]),
    .b(al_fab6b65e[12]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7e1b295f (
    .a(al_c7be2582[26]),
    .b(al_fab6b65e[13]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a32cf9d1 (
    .a(al_c7be2582[27]),
    .b(al_fab6b65e[14]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_47eb555b (
    .a(al_c7be2582[28]),
    .b(al_fab6b65e[15]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_abb726bf (
    .a(al_c7be2582[29]),
    .b(al_fab6b65e[16]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ea1a5ace (
    .a(al_c7be2582[30]),
    .b(al_fab6b65e[17]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_27565bce (
    .a(al_c7be2582[31]),
    .b(al_fab6b65e[18]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bf8379f6 (
    .a(al_c7be2582[32]),
    .b(al_fab6b65e[19]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7084bf6e (
    .a(al_c7be2582[33]),
    .b(al_fab6b65e[20]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3dd74667 (
    .a(al_c7be2582[34]),
    .b(al_fab6b65e[21]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5309dbd3 (
    .a(al_c7be2582[35]),
    .b(al_fab6b65e[22]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_58d193c0 (
    .a(al_c7be2582[36]),
    .b(al_fab6b65e[23]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3a1aeb37 (
    .a(al_c7be2582[37]),
    .b(al_fab6b65e[24]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7d8d958d (
    .a(al_c7be2582[38]),
    .b(al_fab6b65e[25]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9dd45155 (
    .a(al_c7be2582[39]),
    .b(al_fab6b65e[26]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[39]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6a3366e7 (
    .a(al_c7be2582[40]),
    .b(al_fab6b65e[27]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[40]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8551396e (
    .a(al_c7be2582[41]),
    .b(al_fab6b65e[28]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[41]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_414d75a6 (
    .a(al_c7be2582[42]),
    .b(al_fab6b65e[29]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[42]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_97195eda (
    .a(al_c7be2582[43]),
    .b(al_fab6b65e[30]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[43]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1ef82922 (
    .a(al_c7be2582[44]),
    .b(al_fab6b65e[31]),
    .c(al_5b4dd00b),
    .o(al_be68a6d4[44]));
  AL_DFF_X al_62f21365 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[0]));
  AL_DFF_X al_d7b25a44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[9]));
  AL_DFF_X al_1c6460e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[10]));
  AL_DFF_X al_852ecfd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[11]));
  AL_DFF_X al_3235844 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[12]));
  AL_DFF_X al_28335cc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[13]));
  AL_DFF_X al_b015fae1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[14]));
  AL_DFF_X al_b4589968 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[15]));
  AL_DFF_X al_de63bd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[16]));
  AL_DFF_X al_6394b341 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[17]));
  AL_DFF_X al_e0627cd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[18]));
  AL_DFF_X al_90cdf5ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[1]));
  AL_DFF_X al_2df44f6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[19]));
  AL_DFF_X al_b16996a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[20]));
  AL_DFF_X al_46c80a32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[21]));
  AL_DFF_X al_78bcd2ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[22]));
  AL_DFF_X al_194faf5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[23]));
  AL_DFF_X al_8dc74381 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[24]));
  AL_DFF_X al_4d695666 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[25]));
  AL_DFF_X al_e00578bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[26]));
  AL_DFF_X al_5dea13a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[27]));
  AL_DFF_X al_3a3567cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[28]));
  AL_DFF_X al_1a74c879 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[2]));
  AL_DFF_X al_56368394 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[29]));
  AL_DFF_X al_6f220a2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[30]));
  AL_DFF_X al_8fcae728 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[31]));
  AL_DFF_X al_ef257c22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[32]));
  AL_DFF_X al_f2305256 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[33]));
  AL_DFF_X al_74d66024 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[34]));
  AL_DFF_X al_78674213 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[35]));
  AL_DFF_X al_fcbe6479 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[36]));
  AL_DFF_X al_8eb5e728 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[37]));
  AL_DFF_X al_6486f0ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[38]));
  AL_DFF_X al_c7c49285 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[3]));
  AL_DFF_X al_4c16753b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[39]));
  AL_DFF_X al_8fda8ffb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[40]));
  AL_DFF_X al_4c0c28f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[41]));
  AL_DFF_X al_474ecd64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[42]));
  AL_DFF_X al_e48e4e22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[43]));
  AL_DFF_X al_10c26515 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_be68a6d4[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[44]));
  AL_DFF_X al_4ea64755 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[4]));
  AL_DFF_X al_fb0892c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[5]));
  AL_DFF_X al_ba2fab86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[6]));
  AL_DFF_X al_46bcb5f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[7]));
  AL_DFF_X al_ea03efd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c7be2582[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d99b0302[8]));
  AL_DFF_X al_ca203b4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5b4dd00b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[0]));
  AL_DFF_X al_a1b1a461 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[9]));
  AL_DFF_X al_cbf1bfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[10]));
  AL_DFF_X al_b82bd4b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[11]));
  AL_DFF_X al_3f7c497d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[12]));
  AL_DFF_X al_75010a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[13]));
  AL_DFF_X al_69a2cd4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[14]));
  AL_DFF_X al_24a687f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[15]));
  AL_DFF_X al_1ecc244a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[16]));
  AL_DFF_X al_c8fe2b91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[17]));
  AL_DFF_X al_be73cd5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[18]));
  AL_DFF_X al_540f03b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[1]));
  AL_DFF_X al_815f5dbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[19]));
  AL_DFF_X al_40cdac95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[20]));
  AL_DFF_X al_2a1d5196 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[21]));
  AL_DFF_X al_944ac0b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[22]));
  AL_DFF_X al_aa782a7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[23]));
  AL_DFF_X al_33ea299c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[24]));
  AL_DFF_X al_bcbb3972 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[25]));
  AL_DFF_X al_3d81a09c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[26]));
  AL_DFF_X al_16f710c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[27]));
  AL_DFF_X al_f77c792e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[28]));
  AL_DFF_X al_13455c12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[2]));
  AL_DFF_X al_43461d86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[29]));
  AL_DFF_X al_1ba8bcd3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[30]));
  AL_DFF_X al_54d36354 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[31]));
  AL_DFF_X al_7a8d90e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[32]));
  AL_DFF_X al_685fc62f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[33]));
  AL_DFF_X al_42b40ffc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[34]));
  AL_DFF_X al_88f22c71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[3]));
  AL_DFF_X al_14fe75ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[4]));
  AL_DFF_X al_bc0342df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[5]));
  AL_DFF_X al_259b62e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[6]));
  AL_DFF_X al_6a486c91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[7]));
  AL_DFF_X al_3f41cc76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_64e3fb17[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8642d51e[8]));
  AL_DFF_X al_d48ce46a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_65c09044[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4c0a9e6a[0]));
  AL_DFF_X al_742b6587 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[11]));
  AL_DFF_X al_7976e16e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[12]));
  AL_DFF_X al_9f49d72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[13]));
  AL_DFF_X al_3c71ee11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[14]));
  AL_DFF_X al_ed981400 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[15]));
  AL_DFF_X al_81054a97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[16]));
  AL_DFF_X al_9ec4ad5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[17]));
  AL_DFF_X al_98022ea5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[18]));
  AL_DFF_X al_bb184dd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[19]));
  AL_DFF_X al_c0d43797 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[20]));
  AL_DFF_X al_4919f6cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[21]));
  AL_DFF_X al_d37753a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[22]));
  AL_DFF_X al_e8d38d44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[23]));
  AL_DFF_X al_b1de52bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[24]));
  AL_DFF_X al_2395b00f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[25]));
  AL_DFF_X al_9620291c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[26]));
  AL_DFF_X al_158f8b83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[27]));
  AL_DFF_X al_efacaae8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[28]));
  AL_DFF_X al_4338744 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[29]));
  AL_DFF_X al_53a0f96f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[30]));
  AL_DFF_X al_2ec5a207 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[31]));
  AL_DFF_X al_2c17942d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[32]));
  AL_DFF_X al_83e0bae3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[33]));
  AL_DFF_X al_8f885aa3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[34]));
  AL_DFF_X al_1471c412 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[35]));
  AL_DFF_X al_667e5f98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[36]));
  AL_DFF_X al_ccb5432b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[37]));
  AL_DFF_X al_fb673801 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[38]));
  AL_DFF_X al_fe619a17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[39]));
  AL_DFF_X al_26052681 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[40]));
  AL_DFF_X al_b571297f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[41]));
  AL_DFF_X al_2542381a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bac230e2[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ccda870f[42]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_3922abc0 (
    .a(1'b0),
    .o({al_584eea74,open_n147}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3188a5b5 (
    .a(al_d99b0302[12]),
    .b(al_bac230e2[12]),
    .c(al_584eea74),
    .o({al_c6e57848,al_cc14d64d[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ffb0d1f3 (
    .a(al_d99b0302[13]),
    .b(al_bac230e2[13]),
    .c(al_c6e57848),
    .o({al_efc6812a,al_cc14d64d[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_98f6623 (
    .a(al_d99b0302[14]),
    .b(al_bac230e2[14]),
    .c(al_efc6812a),
    .o({al_10825af9,al_cc14d64d[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_26b012e (
    .a(al_d99b0302[15]),
    .b(al_bac230e2[15]),
    .c(al_10825af9),
    .o({al_bbfa0f21,al_cc14d64d[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_369c2d46 (
    .a(al_d99b0302[16]),
    .b(al_bac230e2[16]),
    .c(al_bbfa0f21),
    .o({al_bf9072a4,al_cc14d64d[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_52cbcd99 (
    .a(al_d99b0302[17]),
    .b(al_bac230e2[17]),
    .c(al_bf9072a4),
    .o({al_18cc4352,al_cc14d64d[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_646e468b (
    .a(al_d99b0302[18]),
    .b(al_bac230e2[18]),
    .c(al_18cc4352),
    .o({al_cd59a509,al_cc14d64d[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c68a7283 (
    .a(al_d99b0302[19]),
    .b(al_bac230e2[19]),
    .c(al_cd59a509),
    .o({al_a9bd067e,al_cc14d64d[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d0ecbcb0 (
    .a(al_d99b0302[20]),
    .b(al_bac230e2[20]),
    .c(al_a9bd067e),
    .o({al_8ff81b47,al_cc14d64d[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2c3c2565 (
    .a(al_d99b0302[21]),
    .b(al_bac230e2[21]),
    .c(al_8ff81b47),
    .o({al_91d9bc15,al_cc14d64d[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3dffb78e (
    .a(al_d99b0302[22]),
    .b(al_bac230e2[22]),
    .c(al_91d9bc15),
    .o({al_da758300,al_cc14d64d[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3e2d44eb (
    .a(al_d99b0302[23]),
    .b(al_bac230e2[23]),
    .c(al_da758300),
    .o({al_44b995d2,al_cc14d64d[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c4e0ab9f (
    .a(al_d99b0302[24]),
    .b(al_bac230e2[24]),
    .c(al_44b995d2),
    .o({al_f3c33aa1,al_cc14d64d[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d0e3d41e (
    .a(al_d99b0302[25]),
    .b(al_bac230e2[25]),
    .c(al_f3c33aa1),
    .o({al_1b86bf86,al_cc14d64d[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a24e7f92 (
    .a(al_d99b0302[26]),
    .b(al_bac230e2[26]),
    .c(al_1b86bf86),
    .o({al_d1142aec,al_cc14d64d[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_df013b43 (
    .a(al_d99b0302[27]),
    .b(al_bac230e2[27]),
    .c(al_d1142aec),
    .o({al_6600d0f4,al_cc14d64d[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_aaf1efb2 (
    .a(al_d99b0302[28]),
    .b(al_bac230e2[28]),
    .c(al_6600d0f4),
    .o({al_e73d5abc,al_cc14d64d[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1b618364 (
    .a(al_d99b0302[29]),
    .b(al_bac230e2[29]),
    .c(al_e73d5abc),
    .o({al_a2618249,al_cc14d64d[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_deaf39a6 (
    .a(al_d99b0302[30]),
    .b(al_bac230e2[30]),
    .c(al_a2618249),
    .o({al_e181fe09,al_cc14d64d[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2675a644 (
    .a(al_d99b0302[31]),
    .b(al_bac230e2[31]),
    .c(al_e181fe09),
    .o({al_c77349a0,al_cc14d64d[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dd7547cf (
    .a(al_d99b0302[32]),
    .b(al_bac230e2[32]),
    .c(al_c77349a0),
    .o({al_f63d2d13,al_cc14d64d[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bb326ace (
    .a(al_d99b0302[33]),
    .b(al_bac230e2[33]),
    .c(al_f63d2d13),
    .o({al_46537d2e,al_cc14d64d[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8d037a7a (
    .a(al_d99b0302[34]),
    .b(al_bac230e2[34]),
    .c(al_46537d2e),
    .o({al_a889f4bf,al_cc14d64d[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6c7ba6e (
    .a(al_d99b0302[35]),
    .b(al_bac230e2[35]),
    .c(al_a889f4bf),
    .o({al_accde4d,al_cc14d64d[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9da91bbd (
    .a(al_d99b0302[36]),
    .b(al_bac230e2[36]),
    .c(al_accde4d),
    .o({al_508bf5eb,al_cc14d64d[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2e21c2a6 (
    .a(al_d99b0302[37]),
    .b(al_bac230e2[37]),
    .c(al_508bf5eb),
    .o({al_e82cb205,al_cc14d64d[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_167d0e23 (
    .a(al_d99b0302[38]),
    .b(al_bac230e2[38]),
    .c(al_e82cb205),
    .o({al_4f99c2a2,al_cc14d64d[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e2cb20c (
    .a(al_d99b0302[39]),
    .b(al_bac230e2[39]),
    .c(al_4f99c2a2),
    .o({al_46d116b1,al_cc14d64d[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ebcdf549 (
    .a(al_d99b0302[40]),
    .b(al_bac230e2[40]),
    .c(al_46d116b1),
    .o({al_7a5c8d6e,al_cc14d64d[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_18535c7c (
    .a(al_d99b0302[41]),
    .b(al_bac230e2[41]),
    .c(al_7a5c8d6e),
    .o({al_86d44bba,al_cc14d64d[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d93b520d (
    .a(al_d99b0302[42]),
    .b(al_bac230e2[42]),
    .c(al_86d44bba),
    .o({al_53b3d48f,al_cc14d64d[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e5eedb63 (
    .a(al_d99b0302[43]),
    .b(al_bac230e2[43]),
    .c(al_53b3d48f),
    .o({al_7ed64a67,al_cc14d64d[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1af8a5d5 (
    .a(al_d99b0302[44]),
    .b(1'b0),
    .c(al_7ed64a67),
    .o({al_779d4335,open_n148}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2708e378 (
    .a(1'b0),
    .b(1'b1),
    .c(al_779d4335),
    .o({open_n149,al_e0b2aa1b}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1326908e (
    .a(al_d99b0302[12]),
    .b(al_cc14d64d[0]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_23ed27eb (
    .a(al_d99b0302[13]),
    .b(al_cc14d64d[1]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fd1fa997 (
    .a(al_d99b0302[14]),
    .b(al_cc14d64d[2]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e31c19a9 (
    .a(al_d99b0302[15]),
    .b(al_cc14d64d[3]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1dbe3271 (
    .a(al_d99b0302[16]),
    .b(al_cc14d64d[4]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7f28a8aa (
    .a(al_d99b0302[17]),
    .b(al_cc14d64d[5]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bc27e52c (
    .a(al_d99b0302[18]),
    .b(al_cc14d64d[6]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_57f1b2c (
    .a(al_d99b0302[19]),
    .b(al_cc14d64d[7]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c2103bd6 (
    .a(al_d99b0302[20]),
    .b(al_cc14d64d[8]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_92870231 (
    .a(al_d99b0302[21]),
    .b(al_cc14d64d[9]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3aa59330 (
    .a(al_d99b0302[22]),
    .b(al_cc14d64d[10]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1507efa4 (
    .a(al_d99b0302[23]),
    .b(al_cc14d64d[11]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_12971331 (
    .a(al_d99b0302[24]),
    .b(al_cc14d64d[12]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9a69f626 (
    .a(al_d99b0302[25]),
    .b(al_cc14d64d[13]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b242ca0e (
    .a(al_d99b0302[26]),
    .b(al_cc14d64d[14]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_49e63786 (
    .a(al_d99b0302[27]),
    .b(al_cc14d64d[15]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_172bb920 (
    .a(al_d99b0302[28]),
    .b(al_cc14d64d[16]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7a01e9b9 (
    .a(al_d99b0302[29]),
    .b(al_cc14d64d[17]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f9869f48 (
    .a(al_d99b0302[30]),
    .b(al_cc14d64d[18]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ff210bbb (
    .a(al_d99b0302[31]),
    .b(al_cc14d64d[19]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6644a0d9 (
    .a(al_d99b0302[32]),
    .b(al_cc14d64d[20]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_df63329 (
    .a(al_d99b0302[33]),
    .b(al_cc14d64d[21]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b139b9b5 (
    .a(al_d99b0302[34]),
    .b(al_cc14d64d[22]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ba89dd15 (
    .a(al_d99b0302[35]),
    .b(al_cc14d64d[23]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c8fe4a36 (
    .a(al_d99b0302[36]),
    .b(al_cc14d64d[24]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3530c6b9 (
    .a(al_d99b0302[37]),
    .b(al_cc14d64d[25]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_36cb86a (
    .a(al_d99b0302[38]),
    .b(al_cc14d64d[26]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9b71db1d (
    .a(al_d99b0302[39]),
    .b(al_cc14d64d[27]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[39]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c6b0e3b5 (
    .a(al_d99b0302[40]),
    .b(al_cc14d64d[28]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[40]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_dabc76c3 (
    .a(al_d99b0302[41]),
    .b(al_cc14d64d[29]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[41]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fc683c32 (
    .a(al_d99b0302[42]),
    .b(al_cc14d64d[30]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[42]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2c79886e (
    .a(al_d99b0302[43]),
    .b(al_cc14d64d[31]),
    .c(al_e0b2aa1b),
    .o(al_b75cf8f9[43]));
  AL_DFF_X al_c3c771f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[0]));
  AL_DFF_X al_8501f7aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[9]));
  AL_DFF_X al_8b1a1e0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[10]));
  AL_DFF_X al_ce26601c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[11]));
  AL_DFF_X al_8435049f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[12]));
  AL_DFF_X al_e8573e4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[13]));
  AL_DFF_X al_6411ed1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[14]));
  AL_DFF_X al_4e3223eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[15]));
  AL_DFF_X al_b4712450 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[16]));
  AL_DFF_X al_5e0d236e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[17]));
  AL_DFF_X al_7d56cead (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[18]));
  AL_DFF_X al_83d9dd57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[1]));
  AL_DFF_X al_60db15d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[19]));
  AL_DFF_X al_2567f111 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[20]));
  AL_DFF_X al_bde84bce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[21]));
  AL_DFF_X al_4d7ecfba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[22]));
  AL_DFF_X al_cdce51a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[23]));
  AL_DFF_X al_80c9acd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[24]));
  AL_DFF_X al_ac53a60f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[25]));
  AL_DFF_X al_4c12a30f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[26]));
  AL_DFF_X al_1354590 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[27]));
  AL_DFF_X al_2839745a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[28]));
  AL_DFF_X al_a8c3e901 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[2]));
  AL_DFF_X al_871534fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[29]));
  AL_DFF_X al_49508f5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[30]));
  AL_DFF_X al_d343a789 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[31]));
  AL_DFF_X al_3f535eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[32]));
  AL_DFF_X al_46918f9b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[33]));
  AL_DFF_X al_e9ad6551 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[34]));
  AL_DFF_X al_9804ba4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[35]));
  AL_DFF_X al_c08f1e01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[36]));
  AL_DFF_X al_a623e6df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[37]));
  AL_DFF_X al_3555974f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[38]));
  AL_DFF_X al_33cc389b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[3]));
  AL_DFF_X al_2cd89bf9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[39]));
  AL_DFF_X al_34b748a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[40]));
  AL_DFF_X al_56c25059 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[41]));
  AL_DFF_X al_b9c1325 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[42]));
  AL_DFF_X al_38d2e0f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b75cf8f9[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[43]));
  AL_DFF_X al_e843c648 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[4]));
  AL_DFF_X al_2f99db2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[5]));
  AL_DFF_X al_c0ee3e38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[6]));
  AL_DFF_X al_749c0a05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[7]));
  AL_DFF_X al_a6e55879 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d99b0302[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cb972596[8]));
  AL_DFF_X al_897b894b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e0b2aa1b),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[0]));
  AL_DFF_X al_e8a19370 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[9]));
  AL_DFF_X al_ccb7398 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[10]));
  AL_DFF_X al_3146f4da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[11]));
  AL_DFF_X al_27fe0b4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[12]));
  AL_DFF_X al_fbca34b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[13]));
  AL_DFF_X al_f7c76b5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[14]));
  AL_DFF_X al_8359ce0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[15]));
  AL_DFF_X al_2cd0df1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[16]));
  AL_DFF_X al_fc297270 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[17]));
  AL_DFF_X al_4e567b75 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[18]));
  AL_DFF_X al_a708be8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[1]));
  AL_DFF_X al_82c2e5f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[19]));
  AL_DFF_X al_43fd785b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[20]));
  AL_DFF_X al_5d28a0b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[21]));
  AL_DFF_X al_438de26b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[22]));
  AL_DFF_X al_fc45f2c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[23]));
  AL_DFF_X al_cd1b5918 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[24]));
  AL_DFF_X al_e14f4b65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[25]));
  AL_DFF_X al_fb8de732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[26]));
  AL_DFF_X al_ed2723d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[27]));
  AL_DFF_X al_8fa8a2fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[28]));
  AL_DFF_X al_8c43b4cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[2]));
  AL_DFF_X al_e1745e14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[29]));
  AL_DFF_X al_119fd869 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[30]));
  AL_DFF_X al_46407ab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[31]));
  AL_DFF_X al_6cde6453 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[32]));
  AL_DFF_X al_901b44c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[33]));
  AL_DFF_X al_a2baddea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[34]));
  AL_DFF_X al_1b990587 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[35]));
  AL_DFF_X al_febf1384 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[3]));
  AL_DFF_X al_91d93ee6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[4]));
  AL_DFF_X al_9a420013 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[5]));
  AL_DFF_X al_d5ec03c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[6]));
  AL_DFF_X al_f64404cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[7]));
  AL_DFF_X al_3a9ccbc2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8642d51e[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_29052500[8]));
  AL_DFF_X al_baae8888 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4c0a9e6a[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_88b72b17[0]));
  AL_DFF_X al_d30f614 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[10]));
  AL_DFF_X al_9b6ccacb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[11]));
  AL_DFF_X al_2246f37f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[12]));
  AL_DFF_X al_b677d93e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[13]));
  AL_DFF_X al_383c745f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[14]));
  AL_DFF_X al_3d7901a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[15]));
  AL_DFF_X al_40879df1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[16]));
  AL_DFF_X al_916b01ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[17]));
  AL_DFF_X al_8e2953b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[18]));
  AL_DFF_X al_92cca7af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[19]));
  AL_DFF_X al_2d8bac3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[20]));
  AL_DFF_X al_9dfab16f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[21]));
  AL_DFF_X al_c5e78b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[22]));
  AL_DFF_X al_1f7302d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[23]));
  AL_DFF_X al_b7a2c988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[24]));
  AL_DFF_X al_be802464 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[25]));
  AL_DFF_X al_45900106 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[26]));
  AL_DFF_X al_6de727c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[27]));
  AL_DFF_X al_726e2449 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[28]));
  AL_DFF_X al_9764a957 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[29]));
  AL_DFF_X al_a9f117a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[30]));
  AL_DFF_X al_2f392a8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[31]));
  AL_DFF_X al_e0ade7f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[32]));
  AL_DFF_X al_3be272e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[33]));
  AL_DFF_X al_6f16f2f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[34]));
  AL_DFF_X al_a40bc81b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[35]));
  AL_DFF_X al_a0f6712a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[36]));
  AL_DFF_X al_30851c20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[37]));
  AL_DFF_X al_cc38678f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[38]));
  AL_DFF_X al_d586271e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[39]));
  AL_DFF_X al_7ea44779 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[40]));
  AL_DFF_X al_1171c7ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ccda870f[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8c4c0e00[41]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_92ac89b0 (
    .a(1'b0),
    .o({al_38a13889,open_n152}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9921361f (
    .a(al_cb972596[11]),
    .b(al_ccda870f[11]),
    .c(al_38a13889),
    .o({al_8419f2ed,al_35eab049[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ef3c5115 (
    .a(al_cb972596[12]),
    .b(al_ccda870f[12]),
    .c(al_8419f2ed),
    .o({al_f54b9335,al_35eab049[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8f6ef6e7 (
    .a(al_cb972596[13]),
    .b(al_ccda870f[13]),
    .c(al_f54b9335),
    .o({al_8ed6d91d,al_35eab049[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_def1ef1c (
    .a(al_cb972596[14]),
    .b(al_ccda870f[14]),
    .c(al_8ed6d91d),
    .o({al_3a63fdce,al_35eab049[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e1bebbac (
    .a(al_cb972596[15]),
    .b(al_ccda870f[15]),
    .c(al_3a63fdce),
    .o({al_7d6eed39,al_35eab049[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c05901b2 (
    .a(al_cb972596[16]),
    .b(al_ccda870f[16]),
    .c(al_7d6eed39),
    .o({al_ebfc32c7,al_35eab049[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1398e24b (
    .a(al_cb972596[17]),
    .b(al_ccda870f[17]),
    .c(al_ebfc32c7),
    .o({al_34381ac,al_35eab049[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4ce7182e (
    .a(al_cb972596[18]),
    .b(al_ccda870f[18]),
    .c(al_34381ac),
    .o({al_49175cff,al_35eab049[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_59ecb15d (
    .a(al_cb972596[19]),
    .b(al_ccda870f[19]),
    .c(al_49175cff),
    .o({al_63ff6480,al_35eab049[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ae54cd39 (
    .a(al_cb972596[20]),
    .b(al_ccda870f[20]),
    .c(al_63ff6480),
    .o({al_27dd2411,al_35eab049[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7e9a87a0 (
    .a(al_cb972596[21]),
    .b(al_ccda870f[21]),
    .c(al_27dd2411),
    .o({al_a911db93,al_35eab049[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d0f13c1e (
    .a(al_cb972596[22]),
    .b(al_ccda870f[22]),
    .c(al_a911db93),
    .o({al_405a9f2c,al_35eab049[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_58bc5432 (
    .a(al_cb972596[23]),
    .b(al_ccda870f[23]),
    .c(al_405a9f2c),
    .o({al_e8221400,al_35eab049[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_374990a6 (
    .a(al_cb972596[24]),
    .b(al_ccda870f[24]),
    .c(al_e8221400),
    .o({al_a28a7cde,al_35eab049[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_be60174b (
    .a(al_cb972596[25]),
    .b(al_ccda870f[25]),
    .c(al_a28a7cde),
    .o({al_61046848,al_35eab049[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_32119611 (
    .a(al_cb972596[26]),
    .b(al_ccda870f[26]),
    .c(al_61046848),
    .o({al_51208526,al_35eab049[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9ade1a0e (
    .a(al_cb972596[27]),
    .b(al_ccda870f[27]),
    .c(al_51208526),
    .o({al_93c8ec69,al_35eab049[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_58cf3d96 (
    .a(al_cb972596[28]),
    .b(al_ccda870f[28]),
    .c(al_93c8ec69),
    .o({al_52ebcad4,al_35eab049[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_432b883b (
    .a(al_cb972596[29]),
    .b(al_ccda870f[29]),
    .c(al_52ebcad4),
    .o({al_ed6494a,al_35eab049[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ed00e5cf (
    .a(al_cb972596[30]),
    .b(al_ccda870f[30]),
    .c(al_ed6494a),
    .o({al_7d39bb7d,al_35eab049[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fca53d65 (
    .a(al_cb972596[31]),
    .b(al_ccda870f[31]),
    .c(al_7d39bb7d),
    .o({al_22aeb069,al_35eab049[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e8023cbd (
    .a(al_cb972596[32]),
    .b(al_ccda870f[32]),
    .c(al_22aeb069),
    .o({al_5d314c19,al_35eab049[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_22d5c333 (
    .a(al_cb972596[33]),
    .b(al_ccda870f[33]),
    .c(al_5d314c19),
    .o({al_53a672a,al_35eab049[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_51e4b4c (
    .a(al_cb972596[34]),
    .b(al_ccda870f[34]),
    .c(al_53a672a),
    .o({al_39309161,al_35eab049[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_35027896 (
    .a(al_cb972596[35]),
    .b(al_ccda870f[35]),
    .c(al_39309161),
    .o({al_9a288672,al_35eab049[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_63230116 (
    .a(al_cb972596[36]),
    .b(al_ccda870f[36]),
    .c(al_9a288672),
    .o({al_d2d28755,al_35eab049[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_faf589bd (
    .a(al_cb972596[37]),
    .b(al_ccda870f[37]),
    .c(al_d2d28755),
    .o({al_baeae313,al_35eab049[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ea51b893 (
    .a(al_cb972596[38]),
    .b(al_ccda870f[38]),
    .c(al_baeae313),
    .o({al_63993f05,al_35eab049[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_89bc62a5 (
    .a(al_cb972596[39]),
    .b(al_ccda870f[39]),
    .c(al_63993f05),
    .o({al_b24d98eb,al_35eab049[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fa75ec4b (
    .a(al_cb972596[40]),
    .b(al_ccda870f[40]),
    .c(al_b24d98eb),
    .o({al_89a36400,al_35eab049[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_130658f (
    .a(al_cb972596[41]),
    .b(al_ccda870f[41]),
    .c(al_89a36400),
    .o({al_1a8ff40a,al_35eab049[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5cd1bc44 (
    .a(al_cb972596[42]),
    .b(al_ccda870f[42]),
    .c(al_1a8ff40a),
    .o({al_585d083c,al_35eab049[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c1173245 (
    .a(al_cb972596[43]),
    .b(1'b0),
    .c(al_585d083c),
    .o({al_bada19ee,open_n153}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5bf04055 (
    .a(1'b0),
    .b(1'b1),
    .c(al_bada19ee),
    .o({open_n154,al_3184f1ad}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fdf3d7c7 (
    .a(al_cb972596[11]),
    .b(al_35eab049[0]),
    .c(al_3184f1ad),
    .o(al_dd187023[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c3baecb4 (
    .a(al_cb972596[12]),
    .b(al_35eab049[1]),
    .c(al_3184f1ad),
    .o(al_dd187023[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_95a1bd7b (
    .a(al_cb972596[13]),
    .b(al_35eab049[2]),
    .c(al_3184f1ad),
    .o(al_dd187023[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8591f38b (
    .a(al_cb972596[14]),
    .b(al_35eab049[3]),
    .c(al_3184f1ad),
    .o(al_dd187023[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4aac87d1 (
    .a(al_cb972596[15]),
    .b(al_35eab049[4]),
    .c(al_3184f1ad),
    .o(al_dd187023[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a3402781 (
    .a(al_cb972596[16]),
    .b(al_35eab049[5]),
    .c(al_3184f1ad),
    .o(al_dd187023[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8db0681 (
    .a(al_cb972596[17]),
    .b(al_35eab049[6]),
    .c(al_3184f1ad),
    .o(al_dd187023[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_161ed372 (
    .a(al_cb972596[18]),
    .b(al_35eab049[7]),
    .c(al_3184f1ad),
    .o(al_dd187023[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_41a27fee (
    .a(al_cb972596[19]),
    .b(al_35eab049[8]),
    .c(al_3184f1ad),
    .o(al_dd187023[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_15fad0e (
    .a(al_cb972596[20]),
    .b(al_35eab049[9]),
    .c(al_3184f1ad),
    .o(al_dd187023[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9efc9586 (
    .a(al_cb972596[21]),
    .b(al_35eab049[10]),
    .c(al_3184f1ad),
    .o(al_dd187023[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cb6feedd (
    .a(al_cb972596[22]),
    .b(al_35eab049[11]),
    .c(al_3184f1ad),
    .o(al_dd187023[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_40176de4 (
    .a(al_cb972596[23]),
    .b(al_35eab049[12]),
    .c(al_3184f1ad),
    .o(al_dd187023[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7e51c380 (
    .a(al_cb972596[24]),
    .b(al_35eab049[13]),
    .c(al_3184f1ad),
    .o(al_dd187023[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f536c8c9 (
    .a(al_cb972596[25]),
    .b(al_35eab049[14]),
    .c(al_3184f1ad),
    .o(al_dd187023[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fde35b09 (
    .a(al_cb972596[26]),
    .b(al_35eab049[15]),
    .c(al_3184f1ad),
    .o(al_dd187023[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_167d2ed7 (
    .a(al_cb972596[27]),
    .b(al_35eab049[16]),
    .c(al_3184f1ad),
    .o(al_dd187023[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_90c3092b (
    .a(al_cb972596[28]),
    .b(al_35eab049[17]),
    .c(al_3184f1ad),
    .o(al_dd187023[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f53a5117 (
    .a(al_cb972596[29]),
    .b(al_35eab049[18]),
    .c(al_3184f1ad),
    .o(al_dd187023[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_191a022e (
    .a(al_cb972596[30]),
    .b(al_35eab049[19]),
    .c(al_3184f1ad),
    .o(al_dd187023[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8c55f69b (
    .a(al_cb972596[31]),
    .b(al_35eab049[20]),
    .c(al_3184f1ad),
    .o(al_dd187023[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1489c4a8 (
    .a(al_cb972596[32]),
    .b(al_35eab049[21]),
    .c(al_3184f1ad),
    .o(al_dd187023[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9c97e822 (
    .a(al_cb972596[33]),
    .b(al_35eab049[22]),
    .c(al_3184f1ad),
    .o(al_dd187023[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c1c53d1d (
    .a(al_cb972596[34]),
    .b(al_35eab049[23]),
    .c(al_3184f1ad),
    .o(al_dd187023[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_44f99a92 (
    .a(al_cb972596[35]),
    .b(al_35eab049[24]),
    .c(al_3184f1ad),
    .o(al_dd187023[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_eb504c1 (
    .a(al_cb972596[36]),
    .b(al_35eab049[25]),
    .c(al_3184f1ad),
    .o(al_dd187023[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3e22e763 (
    .a(al_cb972596[37]),
    .b(al_35eab049[26]),
    .c(al_3184f1ad),
    .o(al_dd187023[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b7816c99 (
    .a(al_cb972596[38]),
    .b(al_35eab049[27]),
    .c(al_3184f1ad),
    .o(al_dd187023[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4093dd50 (
    .a(al_cb972596[39]),
    .b(al_35eab049[28]),
    .c(al_3184f1ad),
    .o(al_dd187023[39]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_eeaaa6ca (
    .a(al_cb972596[40]),
    .b(al_35eab049[29]),
    .c(al_3184f1ad),
    .o(al_dd187023[40]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_809b685c (
    .a(al_cb972596[41]),
    .b(al_35eab049[30]),
    .c(al_3184f1ad),
    .o(al_dd187023[41]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8346af08 (
    .a(al_cb972596[42]),
    .b(al_35eab049[31]),
    .c(al_3184f1ad),
    .o(al_dd187023[42]));
  AL_DFF_X al_c1cf6fc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[0]));
  AL_DFF_X al_efe4e0fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[9]));
  AL_DFF_X al_a07930db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[10]));
  AL_DFF_X al_1aa7e7e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[11]));
  AL_DFF_X al_4e2292d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[12]));
  AL_DFF_X al_59b314bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[13]));
  AL_DFF_X al_8b061e26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[14]));
  AL_DFF_X al_eccbfc39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[15]));
  AL_DFF_X al_6fdf009b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[16]));
  AL_DFF_X al_6dc8c03d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[17]));
  AL_DFF_X al_863f0f70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[18]));
  AL_DFF_X al_f6ec121 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[1]));
  AL_DFF_X al_22fb0719 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[19]));
  AL_DFF_X al_f6eb998f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[20]));
  AL_DFF_X al_7fe55d9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[21]));
  AL_DFF_X al_ca0f79be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[22]));
  AL_DFF_X al_fba343c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[23]));
  AL_DFF_X al_4953f266 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[24]));
  AL_DFF_X al_98175929 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[25]));
  AL_DFF_X al_72e079a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[26]));
  AL_DFF_X al_e816dd08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[27]));
  AL_DFF_X al_635efa40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[28]));
  AL_DFF_X al_9ca9d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[2]));
  AL_DFF_X al_e2e201bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[29]));
  AL_DFF_X al_29c0f94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[30]));
  AL_DFF_X al_df637de7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[31]));
  AL_DFF_X al_ab0734bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[32]));
  AL_DFF_X al_6d34df2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[33]));
  AL_DFF_X al_71aa7fce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[34]));
  AL_DFF_X al_35c0f12e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[35]));
  AL_DFF_X al_4dca981a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[36]));
  AL_DFF_X al_23227c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[37]));
  AL_DFF_X al_98d4b19d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[38]));
  AL_DFF_X al_c43c8be3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[3]));
  AL_DFF_X al_c5afdaec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[39]));
  AL_DFF_X al_57792352 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[40]));
  AL_DFF_X al_1cfe16fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[41]));
  AL_DFF_X al_ed4ed5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_dd187023[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[42]));
  AL_DFF_X al_ff94f39c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[4]));
  AL_DFF_X al_82278d78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[5]));
  AL_DFF_X al_8566f5b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[6]));
  AL_DFF_X al_68f5024d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[7]));
  AL_DFF_X al_f9f3487e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cb972596[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7848278f[8]));
  AL_DFF_X al_e1e97d1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3184f1ad),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[0]));
  AL_DFF_X al_18ad43f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[9]));
  AL_DFF_X al_b33f9db3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[10]));
  AL_DFF_X al_742820ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[11]));
  AL_DFF_X al_125b4790 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[12]));
  AL_DFF_X al_de820108 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[13]));
  AL_DFF_X al_fbb74e2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[14]));
  AL_DFF_X al_8a1a7d14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[15]));
  AL_DFF_X al_63b1e3c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[16]));
  AL_DFF_X al_79af27d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[17]));
  AL_DFF_X al_e4e16596 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[18]));
  AL_DFF_X al_35230168 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[1]));
  AL_DFF_X al_770edac0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[19]));
  AL_DFF_X al_ac9d1f8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[20]));
  AL_DFF_X al_c531fac8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[21]));
  AL_DFF_X al_79472495 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[22]));
  AL_DFF_X al_480f5b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[23]));
  AL_DFF_X al_c3941c94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[24]));
  AL_DFF_X al_208313c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[25]));
  AL_DFF_X al_8105ae5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[26]));
  AL_DFF_X al_e9e249ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[27]));
  AL_DFF_X al_cb9d6e6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[28]));
  AL_DFF_X al_da61e6fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[2]));
  AL_DFF_X al_ad227785 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[29]));
  AL_DFF_X al_4eaa999b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[30]));
  AL_DFF_X al_684b5d3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[31]));
  AL_DFF_X al_7684886a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[32]));
  AL_DFF_X al_c7a7b8ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[33]));
  AL_DFF_X al_a5d722de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[34]));
  AL_DFF_X al_1fb7de5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[35]));
  AL_DFF_X al_d5ee4e9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[36]));
  AL_DFF_X al_267d5641 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[3]));
  AL_DFF_X al_798d6d6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[4]));
  AL_DFF_X al_a7ee07a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[5]));
  AL_DFF_X al_2ea9df7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[6]));
  AL_DFF_X al_51468508 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[7]));
  AL_DFF_X al_a6763e57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_29052500[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6cd22c9c[8]));
  AL_DFF_X al_83a9d44d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_88b72b17[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d72cf58c[0]));
  AL_DFF_X al_a32b0d86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[9]));
  AL_DFF_X al_2b70f31d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[10]));
  AL_DFF_X al_7143d47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[11]));
  AL_DFF_X al_6c3f171c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[12]));
  AL_DFF_X al_3df0a904 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[13]));
  AL_DFF_X al_27fff47e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[14]));
  AL_DFF_X al_94abb2b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[15]));
  AL_DFF_X al_a9285152 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[16]));
  AL_DFF_X al_45a805ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[17]));
  AL_DFF_X al_55ce4e60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[18]));
  AL_DFF_X al_8fc9d2a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[19]));
  AL_DFF_X al_7809c7a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[20]));
  AL_DFF_X al_42d8573f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[21]));
  AL_DFF_X al_8378df87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[22]));
  AL_DFF_X al_18060b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[23]));
  AL_DFF_X al_946b0ba9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[24]));
  AL_DFF_X al_34d1e876 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[25]));
  AL_DFF_X al_d0f46ac2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[26]));
  AL_DFF_X al_ebfd5aa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[27]));
  AL_DFF_X al_325daa11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[28]));
  AL_DFF_X al_8b1cf24a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[29]));
  AL_DFF_X al_291bad12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[30]));
  AL_DFF_X al_79722645 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[31]));
  AL_DFF_X al_a93b6b06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[32]));
  AL_DFF_X al_c8007a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[33]));
  AL_DFF_X al_211ece85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[34]));
  AL_DFF_X al_1dfc7fd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[35]));
  AL_DFF_X al_3bdee31c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[36]));
  AL_DFF_X al_3222f03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[37]));
  AL_DFF_X al_ca8bd927 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[38]));
  AL_DFF_X al_91f5e013 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[39]));
  AL_DFF_X al_16d9037a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c4c0e00[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a32146c7[40]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_7b5a4e37 (
    .a(1'b0),
    .o({al_2bfc7bfc,open_n157}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc91a802 (
    .a(al_7848278f[10]),
    .b(al_8c4c0e00[10]),
    .c(al_2bfc7bfc),
    .o({al_e59a7f64,al_c73a14b6[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1d5ec7d7 (
    .a(al_7848278f[11]),
    .b(al_8c4c0e00[11]),
    .c(al_e59a7f64),
    .o({al_5a56dd8c,al_c73a14b6[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2b7013ec (
    .a(al_7848278f[12]),
    .b(al_8c4c0e00[12]),
    .c(al_5a56dd8c),
    .o({al_c8cc3a74,al_c73a14b6[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1687ffde (
    .a(al_7848278f[13]),
    .b(al_8c4c0e00[13]),
    .c(al_c8cc3a74),
    .o({al_2a0ec313,al_c73a14b6[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_66acd425 (
    .a(al_7848278f[14]),
    .b(al_8c4c0e00[14]),
    .c(al_2a0ec313),
    .o({al_e6e3c466,al_c73a14b6[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5c05c757 (
    .a(al_7848278f[15]),
    .b(al_8c4c0e00[15]),
    .c(al_e6e3c466),
    .o({al_d781087a,al_c73a14b6[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f7aac6e7 (
    .a(al_7848278f[16]),
    .b(al_8c4c0e00[16]),
    .c(al_d781087a),
    .o({al_8cba2b5a,al_c73a14b6[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6d43164 (
    .a(al_7848278f[17]),
    .b(al_8c4c0e00[17]),
    .c(al_8cba2b5a),
    .o({al_cb8ad3a1,al_c73a14b6[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_84fb9a7f (
    .a(al_7848278f[18]),
    .b(al_8c4c0e00[18]),
    .c(al_cb8ad3a1),
    .o({al_3c5da63,al_c73a14b6[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ec981462 (
    .a(al_7848278f[19]),
    .b(al_8c4c0e00[19]),
    .c(al_3c5da63),
    .o({al_731d9b96,al_c73a14b6[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_85fb3344 (
    .a(al_7848278f[20]),
    .b(al_8c4c0e00[20]),
    .c(al_731d9b96),
    .o({al_bf6ae1e2,al_c73a14b6[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_66a1fecc (
    .a(al_7848278f[21]),
    .b(al_8c4c0e00[21]),
    .c(al_bf6ae1e2),
    .o({al_714663e5,al_c73a14b6[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_12c109f6 (
    .a(al_7848278f[22]),
    .b(al_8c4c0e00[22]),
    .c(al_714663e5),
    .o({al_4cf28725,al_c73a14b6[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_41746262 (
    .a(al_7848278f[23]),
    .b(al_8c4c0e00[23]),
    .c(al_4cf28725),
    .o({al_639c27a1,al_c73a14b6[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c0513336 (
    .a(al_7848278f[24]),
    .b(al_8c4c0e00[24]),
    .c(al_639c27a1),
    .o({al_c465640a,al_c73a14b6[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2869e030 (
    .a(al_7848278f[25]),
    .b(al_8c4c0e00[25]),
    .c(al_c465640a),
    .o({al_d013c2db,al_c73a14b6[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1900d99b (
    .a(al_7848278f[26]),
    .b(al_8c4c0e00[26]),
    .c(al_d013c2db),
    .o({al_86c1a1f7,al_c73a14b6[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1f156575 (
    .a(al_7848278f[27]),
    .b(al_8c4c0e00[27]),
    .c(al_86c1a1f7),
    .o({al_e412eb65,al_c73a14b6[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_50f204be (
    .a(al_7848278f[28]),
    .b(al_8c4c0e00[28]),
    .c(al_e412eb65),
    .o({al_f01a65dd,al_c73a14b6[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bcf998bc (
    .a(al_7848278f[29]),
    .b(al_8c4c0e00[29]),
    .c(al_f01a65dd),
    .o({al_e6ba2112,al_c73a14b6[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1825d927 (
    .a(al_7848278f[30]),
    .b(al_8c4c0e00[30]),
    .c(al_e6ba2112),
    .o({al_3fdd05cb,al_c73a14b6[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67569616 (
    .a(al_7848278f[31]),
    .b(al_8c4c0e00[31]),
    .c(al_3fdd05cb),
    .o({al_43bdc053,al_c73a14b6[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_131ee9e5 (
    .a(al_7848278f[32]),
    .b(al_8c4c0e00[32]),
    .c(al_43bdc053),
    .o({al_be037ee1,al_c73a14b6[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_697dddb0 (
    .a(al_7848278f[33]),
    .b(al_8c4c0e00[33]),
    .c(al_be037ee1),
    .o({al_e6e34f55,al_c73a14b6[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_92fd3e23 (
    .a(al_7848278f[34]),
    .b(al_8c4c0e00[34]),
    .c(al_e6e34f55),
    .o({al_a638954c,al_c73a14b6[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4c9fb54 (
    .a(al_7848278f[35]),
    .b(al_8c4c0e00[35]),
    .c(al_a638954c),
    .o({al_9eeedd82,al_c73a14b6[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_409be4d5 (
    .a(al_7848278f[36]),
    .b(al_8c4c0e00[36]),
    .c(al_9eeedd82),
    .o({al_58c037cd,al_c73a14b6[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6aa90d3f (
    .a(al_7848278f[37]),
    .b(al_8c4c0e00[37]),
    .c(al_58c037cd),
    .o({al_f841ecaa,al_c73a14b6[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d5cd0b6f (
    .a(al_7848278f[38]),
    .b(al_8c4c0e00[38]),
    .c(al_f841ecaa),
    .o({al_e7643d65,al_c73a14b6[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ccf35c2a (
    .a(al_7848278f[39]),
    .b(al_8c4c0e00[39]),
    .c(al_e7643d65),
    .o({al_d681bdcc,al_c73a14b6[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_53306aa2 (
    .a(al_7848278f[40]),
    .b(al_8c4c0e00[40]),
    .c(al_d681bdcc),
    .o({al_537d0180,al_c73a14b6[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_42785643 (
    .a(al_7848278f[41]),
    .b(al_8c4c0e00[41]),
    .c(al_537d0180),
    .o({al_c18839e1,al_c73a14b6[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_81a8eacf (
    .a(al_7848278f[42]),
    .b(1'b0),
    .c(al_c18839e1),
    .o({al_a12bfe23,open_n158}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d8df823d (
    .a(1'b0),
    .b(1'b1),
    .c(al_a12bfe23),
    .o({open_n159,al_23bcebc4}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9e9955b (
    .a(al_7848278f[10]),
    .b(al_c73a14b6[0]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_371364a5 (
    .a(al_7848278f[11]),
    .b(al_c73a14b6[1]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4f9af469 (
    .a(al_7848278f[12]),
    .b(al_c73a14b6[2]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d3ed9df9 (
    .a(al_7848278f[13]),
    .b(al_c73a14b6[3]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cf941448 (
    .a(al_7848278f[14]),
    .b(al_c73a14b6[4]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4cc0c4dc (
    .a(al_7848278f[15]),
    .b(al_c73a14b6[5]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_49896960 (
    .a(al_7848278f[16]),
    .b(al_c73a14b6[6]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_22d62959 (
    .a(al_7848278f[17]),
    .b(al_c73a14b6[7]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4019b6d1 (
    .a(al_7848278f[18]),
    .b(al_c73a14b6[8]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c9a5fcea (
    .a(al_7848278f[19]),
    .b(al_c73a14b6[9]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c2c2af52 (
    .a(al_7848278f[20]),
    .b(al_c73a14b6[10]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_63e9c4c7 (
    .a(al_7848278f[21]),
    .b(al_c73a14b6[11]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3bfeb6af (
    .a(al_7848278f[22]),
    .b(al_c73a14b6[12]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1daac10a (
    .a(al_7848278f[23]),
    .b(al_c73a14b6[13]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_19f1017a (
    .a(al_7848278f[24]),
    .b(al_c73a14b6[14]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c884e80 (
    .a(al_7848278f[25]),
    .b(al_c73a14b6[15]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_57132aee (
    .a(al_7848278f[26]),
    .b(al_c73a14b6[16]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_61f54be0 (
    .a(al_7848278f[27]),
    .b(al_c73a14b6[17]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a84d956c (
    .a(al_7848278f[28]),
    .b(al_c73a14b6[18]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_de7f7e1a (
    .a(al_7848278f[29]),
    .b(al_c73a14b6[19]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d15c7837 (
    .a(al_7848278f[30]),
    .b(al_c73a14b6[20]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9eb9585 (
    .a(al_7848278f[31]),
    .b(al_c73a14b6[21]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5a4f6f8a (
    .a(al_7848278f[32]),
    .b(al_c73a14b6[22]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d1024069 (
    .a(al_7848278f[33]),
    .b(al_c73a14b6[23]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_779a55bc (
    .a(al_7848278f[34]),
    .b(al_c73a14b6[24]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_73046ee2 (
    .a(al_7848278f[35]),
    .b(al_c73a14b6[25]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d77a629e (
    .a(al_7848278f[36]),
    .b(al_c73a14b6[26]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4d1a4f0e (
    .a(al_7848278f[37]),
    .b(al_c73a14b6[27]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a246130b (
    .a(al_7848278f[38]),
    .b(al_c73a14b6[28]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9ec9ffe1 (
    .a(al_7848278f[39]),
    .b(al_c73a14b6[29]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[39]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_501670d3 (
    .a(al_7848278f[40]),
    .b(al_c73a14b6[30]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[40]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5f9eac6e (
    .a(al_7848278f[41]),
    .b(al_c73a14b6[31]),
    .c(al_23bcebc4),
    .o(al_b8e7a164[41]));
  AL_DFF_X al_27110919 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[0]));
  AL_DFF_X al_2251f831 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[9]));
  AL_DFF_X al_7dc50fb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[10]));
  AL_DFF_X al_37fd4290 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[11]));
  AL_DFF_X al_3d608492 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[12]));
  AL_DFF_X al_635461f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[13]));
  AL_DFF_X al_82ec55db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[14]));
  AL_DFF_X al_f355d809 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[15]));
  AL_DFF_X al_96334a21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[16]));
  AL_DFF_X al_5c497650 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[17]));
  AL_DFF_X al_7b63043d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[18]));
  AL_DFF_X al_34ffc4b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[1]));
  AL_DFF_X al_ed7626e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[19]));
  AL_DFF_X al_b01e79ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[20]));
  AL_DFF_X al_c93c6d78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[21]));
  AL_DFF_X al_ebb98a07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[22]));
  AL_DFF_X al_32326785 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[23]));
  AL_DFF_X al_34ef7e33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[24]));
  AL_DFF_X al_8a35a45c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[25]));
  AL_DFF_X al_4e785f05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[26]));
  AL_DFF_X al_e4e5b934 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[27]));
  AL_DFF_X al_3905006 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[28]));
  AL_DFF_X al_73938a6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[2]));
  AL_DFF_X al_1c1b8ca6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[29]));
  AL_DFF_X al_a228aec6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[30]));
  AL_DFF_X al_8d137514 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[31]));
  AL_DFF_X al_700e10cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[32]));
  AL_DFF_X al_5ad5f5d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[33]));
  AL_DFF_X al_ac6fba05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[34]));
  AL_DFF_X al_bce7d040 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[35]));
  AL_DFF_X al_d4cfd270 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[36]));
  AL_DFF_X al_73e4ccae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[37]));
  AL_DFF_X al_750556f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[38]));
  AL_DFF_X al_4fc70dc3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[3]));
  AL_DFF_X al_10de0bfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[39]));
  AL_DFF_X al_7d9d46eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[40]));
  AL_DFF_X al_9127edc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b8e7a164[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[41]));
  AL_DFF_X al_9f2a11d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[4]));
  AL_DFF_X al_42043361 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[5]));
  AL_DFF_X al_dce17ee1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[6]));
  AL_DFF_X al_21a74cbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[7]));
  AL_DFF_X al_8d21e7bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7848278f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ab78d0a0[8]));
  AL_DFF_X al_6863cd34 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_23bcebc4),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[0]));
  AL_DFF_X al_e5a02b51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[9]));
  AL_DFF_X al_39655c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[10]));
  AL_DFF_X al_7155d105 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[11]));
  AL_DFF_X al_f88fcad7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[12]));
  AL_DFF_X al_160934b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[13]));
  AL_DFF_X al_65555332 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[14]));
  AL_DFF_X al_ce4c5732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[15]));
  AL_DFF_X al_58327525 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[16]));
  AL_DFF_X al_d9760827 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[17]));
  AL_DFF_X al_518faa14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[18]));
  AL_DFF_X al_c4557e69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[1]));
  AL_DFF_X al_6361f8c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[19]));
  AL_DFF_X al_736bb2f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[20]));
  AL_DFF_X al_2d421100 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[21]));
  AL_DFF_X al_9b393b95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[22]));
  AL_DFF_X al_e9bed325 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[23]));
  AL_DFF_X al_3d958a24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[24]));
  AL_DFF_X al_9ca35887 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[25]));
  AL_DFF_X al_4c56951b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[26]));
  AL_DFF_X al_91ff705d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[27]));
  AL_DFF_X al_be91aeb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[28]));
  AL_DFF_X al_9eaef95d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[2]));
  AL_DFF_X al_a5cf866e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[29]));
  AL_DFF_X al_a472051 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[30]));
  AL_DFF_X al_a3acfdcd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[31]));
  AL_DFF_X al_dfab792d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[32]));
  AL_DFF_X al_8aa2b723 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[33]));
  AL_DFF_X al_90fdf0bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[34]));
  AL_DFF_X al_9c447751 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[35]));
  AL_DFF_X al_38f9729d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[36]));
  AL_DFF_X al_cffd0729 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[37]));
  AL_DFF_X al_7c8bad3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[3]));
  AL_DFF_X al_10c0d97b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[4]));
  AL_DFF_X al_81295d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[5]));
  AL_DFF_X al_6a904d48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[6]));
  AL_DFF_X al_db75b782 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[7]));
  AL_DFF_X al_90778732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cd22c9c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5dd36af2[8]));
  AL_DFF_X al_cfb0ed49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d72cf58c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_90e1f6ef[0]));
  AL_DFF_X al_99b80607 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[9]));
  AL_DFF_X al_7fac2c50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[10]));
  AL_DFF_X al_4633e24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[11]));
  AL_DFF_X al_93f7e05d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[12]));
  AL_DFF_X al_99a723ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[13]));
  AL_DFF_X al_13dbb28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[14]));
  AL_DFF_X al_3d2b85a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[15]));
  AL_DFF_X al_2baad6ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[16]));
  AL_DFF_X al_e9a81d68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[17]));
  AL_DFF_X al_a28fcbfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[18]));
  AL_DFF_X al_68c21ce9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[19]));
  AL_DFF_X al_7756e779 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[20]));
  AL_DFF_X al_8264e1a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[21]));
  AL_DFF_X al_6f0b476e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[22]));
  AL_DFF_X al_fbdef08f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[23]));
  AL_DFF_X al_4d909128 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[24]));
  AL_DFF_X al_9116bcf1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[25]));
  AL_DFF_X al_727c670d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[26]));
  AL_DFF_X al_1cd0f65b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[27]));
  AL_DFF_X al_cfcca1f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[28]));
  AL_DFF_X al_1767834e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[29]));
  AL_DFF_X al_3bc5cd1b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[30]));
  AL_DFF_X al_8966463b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[31]));
  AL_DFF_X al_c60b9eb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[32]));
  AL_DFF_X al_d80959d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[33]));
  AL_DFF_X al_337b7e2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[34]));
  AL_DFF_X al_17bb9edf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[35]));
  AL_DFF_X al_2be6ad97 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[36]));
  AL_DFF_X al_d2ed43d2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[37]));
  AL_DFF_X al_6cf30158 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[38]));
  AL_DFF_X al_20ce945d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[39]));
  AL_DFF_X al_d7a18ed1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a32146c7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2ecc3265[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_ae41c043 (
    .a(1'b0),
    .o({al_94fa0ad9,open_n162}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d712ba20 (
    .a(al_ab78d0a0[9]),
    .b(al_a32146c7[9]),
    .c(al_94fa0ad9),
    .o({al_3773fc04,al_d4021fa0[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8a1db398 (
    .a(al_ab78d0a0[10]),
    .b(al_a32146c7[10]),
    .c(al_3773fc04),
    .o({al_8eedc273,al_d4021fa0[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fbb3275f (
    .a(al_ab78d0a0[11]),
    .b(al_a32146c7[11]),
    .c(al_8eedc273),
    .o({al_bd0a1f9d,al_d4021fa0[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_627df433 (
    .a(al_ab78d0a0[12]),
    .b(al_a32146c7[12]),
    .c(al_bd0a1f9d),
    .o({al_48931d43,al_d4021fa0[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b0450c1b (
    .a(al_ab78d0a0[13]),
    .b(al_a32146c7[13]),
    .c(al_48931d43),
    .o({al_bc9b0eaa,al_d4021fa0[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_48a20f09 (
    .a(al_ab78d0a0[14]),
    .b(al_a32146c7[14]),
    .c(al_bc9b0eaa),
    .o({al_35d02980,al_d4021fa0[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_55a281db (
    .a(al_ab78d0a0[15]),
    .b(al_a32146c7[15]),
    .c(al_35d02980),
    .o({al_fee10e00,al_d4021fa0[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f9b1328d (
    .a(al_ab78d0a0[16]),
    .b(al_a32146c7[16]),
    .c(al_fee10e00),
    .o({al_56671d76,al_d4021fa0[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bd03ef2a (
    .a(al_ab78d0a0[17]),
    .b(al_a32146c7[17]),
    .c(al_56671d76),
    .o({al_912d325d,al_d4021fa0[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f2879e27 (
    .a(al_ab78d0a0[18]),
    .b(al_a32146c7[18]),
    .c(al_912d325d),
    .o({al_9f5bba13,al_d4021fa0[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4ae4392d (
    .a(al_ab78d0a0[19]),
    .b(al_a32146c7[19]),
    .c(al_9f5bba13),
    .o({al_93b8640e,al_d4021fa0[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c9d5405e (
    .a(al_ab78d0a0[20]),
    .b(al_a32146c7[20]),
    .c(al_93b8640e),
    .o({al_e3447775,al_d4021fa0[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_da4a6893 (
    .a(al_ab78d0a0[21]),
    .b(al_a32146c7[21]),
    .c(al_e3447775),
    .o({al_ba94a953,al_d4021fa0[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d462d6b (
    .a(al_ab78d0a0[22]),
    .b(al_a32146c7[22]),
    .c(al_ba94a953),
    .o({al_75a96ab5,al_d4021fa0[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6f0a7e12 (
    .a(al_ab78d0a0[23]),
    .b(al_a32146c7[23]),
    .c(al_75a96ab5),
    .o({al_3c16a30a,al_d4021fa0[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e9ddc85d (
    .a(al_ab78d0a0[24]),
    .b(al_a32146c7[24]),
    .c(al_3c16a30a),
    .o({al_fdf3ddc7,al_d4021fa0[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_be9d8bfe (
    .a(al_ab78d0a0[25]),
    .b(al_a32146c7[25]),
    .c(al_fdf3ddc7),
    .o({al_2c40a92e,al_d4021fa0[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_46152546 (
    .a(al_ab78d0a0[26]),
    .b(al_a32146c7[26]),
    .c(al_2c40a92e),
    .o({al_d57289de,al_d4021fa0[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e166b2f (
    .a(al_ab78d0a0[27]),
    .b(al_a32146c7[27]),
    .c(al_d57289de),
    .o({al_c0464485,al_d4021fa0[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1d1cb04a (
    .a(al_ab78d0a0[28]),
    .b(al_a32146c7[28]),
    .c(al_c0464485),
    .o({al_6cd1bb56,al_d4021fa0[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e098951f (
    .a(al_ab78d0a0[29]),
    .b(al_a32146c7[29]),
    .c(al_6cd1bb56),
    .o({al_805eafcd,al_d4021fa0[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a9284b3 (
    .a(al_ab78d0a0[30]),
    .b(al_a32146c7[30]),
    .c(al_805eafcd),
    .o({al_afc2f09b,al_d4021fa0[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d2fb04e5 (
    .a(al_ab78d0a0[31]),
    .b(al_a32146c7[31]),
    .c(al_afc2f09b),
    .o({al_b626be09,al_d4021fa0[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8ef40365 (
    .a(al_ab78d0a0[32]),
    .b(al_a32146c7[32]),
    .c(al_b626be09),
    .o({al_47857556,al_d4021fa0[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_25d8b345 (
    .a(al_ab78d0a0[33]),
    .b(al_a32146c7[33]),
    .c(al_47857556),
    .o({al_cdf5386d,al_d4021fa0[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_35259b8f (
    .a(al_ab78d0a0[34]),
    .b(al_a32146c7[34]),
    .c(al_cdf5386d),
    .o({al_44a63fb7,al_d4021fa0[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4386b6b0 (
    .a(al_ab78d0a0[35]),
    .b(al_a32146c7[35]),
    .c(al_44a63fb7),
    .o({al_d8fe84e6,al_d4021fa0[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7917d94f (
    .a(al_ab78d0a0[36]),
    .b(al_a32146c7[36]),
    .c(al_d8fe84e6),
    .o({al_6d9bce46,al_d4021fa0[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eddfce27 (
    .a(al_ab78d0a0[37]),
    .b(al_a32146c7[37]),
    .c(al_6d9bce46),
    .o({al_46c8a269,al_d4021fa0[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_168bd9cb (
    .a(al_ab78d0a0[38]),
    .b(al_a32146c7[38]),
    .c(al_46c8a269),
    .o({al_ba4595c0,al_d4021fa0[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a31b4798 (
    .a(al_ab78d0a0[39]),
    .b(al_a32146c7[39]),
    .c(al_ba4595c0),
    .o({al_5bf37252,al_d4021fa0[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5df7c8aa (
    .a(al_ab78d0a0[40]),
    .b(al_a32146c7[40]),
    .c(al_5bf37252),
    .o({al_8cb44011,al_d4021fa0[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bf059000 (
    .a(al_ab78d0a0[41]),
    .b(1'b0),
    .c(al_8cb44011),
    .o({al_b5df3e43,open_n163}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_72b4610a (
    .a(1'b0),
    .b(1'b1),
    .c(al_b5df3e43),
    .o({open_n164,al_2392f558}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_62a02958 (
    .a(al_ab78d0a0[10]),
    .b(al_d4021fa0[1]),
    .c(al_2392f558),
    .o(al_1dac5d46[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1bbcf345 (
    .a(al_ab78d0a0[11]),
    .b(al_d4021fa0[2]),
    .c(al_2392f558),
    .o(al_1dac5d46[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bde05635 (
    .a(al_ab78d0a0[12]),
    .b(al_d4021fa0[3]),
    .c(al_2392f558),
    .o(al_1dac5d46[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f488ce33 (
    .a(al_ab78d0a0[13]),
    .b(al_d4021fa0[4]),
    .c(al_2392f558),
    .o(al_1dac5d46[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4ab8973e (
    .a(al_ab78d0a0[14]),
    .b(al_d4021fa0[5]),
    .c(al_2392f558),
    .o(al_1dac5d46[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3f05340f (
    .a(al_ab78d0a0[15]),
    .b(al_d4021fa0[6]),
    .c(al_2392f558),
    .o(al_1dac5d46[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ae7306c8 (
    .a(al_ab78d0a0[16]),
    .b(al_d4021fa0[7]),
    .c(al_2392f558),
    .o(al_1dac5d46[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6417865b (
    .a(al_ab78d0a0[17]),
    .b(al_d4021fa0[8]),
    .c(al_2392f558),
    .o(al_1dac5d46[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fe66dbaf (
    .a(al_ab78d0a0[18]),
    .b(al_d4021fa0[9]),
    .c(al_2392f558),
    .o(al_1dac5d46[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fb27bc2e (
    .a(al_ab78d0a0[19]),
    .b(al_d4021fa0[10]),
    .c(al_2392f558),
    .o(al_1dac5d46[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_878b3300 (
    .a(al_ab78d0a0[20]),
    .b(al_d4021fa0[11]),
    .c(al_2392f558),
    .o(al_1dac5d46[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a7b6cacc (
    .a(al_ab78d0a0[21]),
    .b(al_d4021fa0[12]),
    .c(al_2392f558),
    .o(al_1dac5d46[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5f3968d1 (
    .a(al_ab78d0a0[22]),
    .b(al_d4021fa0[13]),
    .c(al_2392f558),
    .o(al_1dac5d46[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_56ec608e (
    .a(al_ab78d0a0[23]),
    .b(al_d4021fa0[14]),
    .c(al_2392f558),
    .o(al_1dac5d46[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f9ace108 (
    .a(al_ab78d0a0[24]),
    .b(al_d4021fa0[15]),
    .c(al_2392f558),
    .o(al_1dac5d46[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7765223d (
    .a(al_ab78d0a0[25]),
    .b(al_d4021fa0[16]),
    .c(al_2392f558),
    .o(al_1dac5d46[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_914d307f (
    .a(al_ab78d0a0[26]),
    .b(al_d4021fa0[17]),
    .c(al_2392f558),
    .o(al_1dac5d46[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ec6a0b90 (
    .a(al_ab78d0a0[27]),
    .b(al_d4021fa0[18]),
    .c(al_2392f558),
    .o(al_1dac5d46[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_157ee61 (
    .a(al_ab78d0a0[28]),
    .b(al_d4021fa0[19]),
    .c(al_2392f558),
    .o(al_1dac5d46[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5899298 (
    .a(al_ab78d0a0[29]),
    .b(al_d4021fa0[20]),
    .c(al_2392f558),
    .o(al_1dac5d46[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ae26dd5d (
    .a(al_ab78d0a0[30]),
    .b(al_d4021fa0[21]),
    .c(al_2392f558),
    .o(al_1dac5d46[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d320c9e6 (
    .a(al_ab78d0a0[31]),
    .b(al_d4021fa0[22]),
    .c(al_2392f558),
    .o(al_1dac5d46[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_502798e2 (
    .a(al_ab78d0a0[32]),
    .b(al_d4021fa0[23]),
    .c(al_2392f558),
    .o(al_1dac5d46[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4cc1e5f1 (
    .a(al_ab78d0a0[33]),
    .b(al_d4021fa0[24]),
    .c(al_2392f558),
    .o(al_1dac5d46[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8437e30 (
    .a(al_ab78d0a0[34]),
    .b(al_d4021fa0[25]),
    .c(al_2392f558),
    .o(al_1dac5d46[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7febfd0 (
    .a(al_ab78d0a0[35]),
    .b(al_d4021fa0[26]),
    .c(al_2392f558),
    .o(al_1dac5d46[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6cb1849b (
    .a(al_ab78d0a0[36]),
    .b(al_d4021fa0[27]),
    .c(al_2392f558),
    .o(al_1dac5d46[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cb07aed1 (
    .a(al_ab78d0a0[37]),
    .b(al_d4021fa0[28]),
    .c(al_2392f558),
    .o(al_1dac5d46[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_43845f2e (
    .a(al_ab78d0a0[38]),
    .b(al_d4021fa0[29]),
    .c(al_2392f558),
    .o(al_1dac5d46[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_60160bd4 (
    .a(al_ab78d0a0[39]),
    .b(al_d4021fa0[30]),
    .c(al_2392f558),
    .o(al_1dac5d46[39]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7866e1af (
    .a(al_ab78d0a0[40]),
    .b(al_d4021fa0[31]),
    .c(al_2392f558),
    .o(al_1dac5d46[40]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_aaceb475 (
    .a(al_ab78d0a0[9]),
    .b(al_d4021fa0[0]),
    .c(al_2392f558),
    .o(al_1dac5d46[9]));
  AL_DFF_X al_994b3b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ab78d0a0[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[0]));
  AL_DFF_X al_f50aed44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[9]));
  AL_DFF_X al_dc65df0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[10]));
  AL_DFF_X al_7dc51921 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[11]));
  AL_DFF_X al_b189b582 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[12]));
  AL_DFF_X al_104bdf78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[13]));
  AL_DFF_X al_13d2842e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[14]));
  AL_DFF_X al_942b8382 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[15]));
  AL_DFF_X al_24d8446e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[16]));
  AL_DFF_X al_63fb28ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[17]));
  AL_DFF_X al_2238d337 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[18]));
  AL_DFF_X al_41a1b5c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ab78d0a0[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[1]));
  AL_DFF_X al_fc58b64f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[19]));
  AL_DFF_X al_ba5ed016 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[20]));
  AL_DFF_X al_a0060ca7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[21]));
  AL_DFF_X al_cc027f3f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[22]));
  AL_DFF_X al_63510ff9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[23]));
  AL_DFF_X al_258af1f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[24]));
  AL_DFF_X al_1de87f57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[25]));
  AL_DFF_X al_279ecd26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[26]));
  AL_DFF_X al_4d420542 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[27]));
  AL_DFF_X al_5ceabc3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[28]));
  AL_DFF_X al_c7ceb617 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ab78d0a0[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[2]));
  AL_DFF_X al_fa7c9436 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[29]));
  AL_DFF_X al_f5055da3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[30]));
  AL_DFF_X al_409aebd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[31]));
  AL_DFF_X al_2e0f8d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[32]));
  AL_DFF_X al_7b816eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[33]));
  AL_DFF_X al_a7427e01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[34]));
  AL_DFF_X al_a42ee3c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[35]));
  AL_DFF_X al_48b4c988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[36]));
  AL_DFF_X al_f54e77dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[37]));
  AL_DFF_X al_de8aed86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[38]));
  AL_DFF_X al_85fe55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ab78d0a0[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[3]));
  AL_DFF_X al_31a460a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[39]));
  AL_DFF_X al_bc06f5c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1dac5d46[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[40]));
  AL_DFF_X al_f2eb6f84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ab78d0a0[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[4]));
  AL_DFF_X al_22014898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ab78d0a0[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[5]));
  AL_DFF_X al_d77bc416 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ab78d0a0[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[6]));
  AL_DFF_X al_a3c4056b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ab78d0a0[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[7]));
  AL_DFF_X al_715ca214 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ab78d0a0[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7af0d249[8]));
  AL_DFF_X al_52b73370 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2392f558),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[0]));
  AL_DFF_X al_16de7173 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[9]));
  AL_DFF_X al_78c3857d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[10]));
  AL_DFF_X al_90cfd43a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[11]));
  AL_DFF_X al_7c2308f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[12]));
  AL_DFF_X al_7ee8403d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[13]));
  AL_DFF_X al_2f12ad13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[14]));
  AL_DFF_X al_b9c064c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[15]));
  AL_DFF_X al_6aa2fad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[16]));
  AL_DFF_X al_86aed3df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[17]));
  AL_DFF_X al_293eed6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[18]));
  AL_DFF_X al_c6fe9c43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[1]));
  AL_DFF_X al_863df23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[19]));
  AL_DFF_X al_66ab0e52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[20]));
  AL_DFF_X al_c3ecc727 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[21]));
  AL_DFF_X al_9b1d4969 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[22]));
  AL_DFF_X al_5e17ffc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[23]));
  AL_DFF_X al_5ed1e49a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[24]));
  AL_DFF_X al_1911c075 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[25]));
  AL_DFF_X al_5fbf4b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[26]));
  AL_DFF_X al_682223ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[27]));
  AL_DFF_X al_731138f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[28]));
  AL_DFF_X al_639e5a92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[2]));
  AL_DFF_X al_88b9c53e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[29]));
  AL_DFF_X al_492a9417 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[30]));
  AL_DFF_X al_892693ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[31]));
  AL_DFF_X al_99f1a8ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[32]));
  AL_DFF_X al_fd626b35 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[33]));
  AL_DFF_X al_bbb6c80f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[34]));
  AL_DFF_X al_2d1c7dfd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[35]));
  AL_DFF_X al_3a83de1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[36]));
  AL_DFF_X al_2e5b2bda (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[37]));
  AL_DFF_X al_d0d9e1bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[38]));
  AL_DFF_X al_9816bd1f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[3]));
  AL_DFF_X al_b3eb39a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[4]));
  AL_DFF_X al_3f6a4aa0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[5]));
  AL_DFF_X al_4c64da74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[6]));
  AL_DFF_X al_e6b60508 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[7]));
  AL_DFF_X al_29efc1ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dd36af2[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_b6775e93[8]));
  AL_DFF_X al_5a2d9cf0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_90e1f6ef[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5bcbf559[0]));
  AL_DFF_X al_49825612 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[9]));
  AL_DFF_X al_ad62c7a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[10]));
  AL_DFF_X al_9b18e319 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[11]));
  AL_DFF_X al_ce586cb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[12]));
  AL_DFF_X al_d0d1fa40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[13]));
  AL_DFF_X al_473d1765 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[14]));
  AL_DFF_X al_6bf149e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[15]));
  AL_DFF_X al_879edc39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[16]));
  AL_DFF_X al_d1cc6097 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[17]));
  AL_DFF_X al_bedb2741 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[18]));
  AL_DFF_X al_dfbf5974 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[19]));
  AL_DFF_X al_827ad742 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[20]));
  AL_DFF_X al_9f879568 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[21]));
  AL_DFF_X al_a3fa476f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[22]));
  AL_DFF_X al_513303fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[23]));
  AL_DFF_X al_ebfe1334 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[24]));
  AL_DFF_X al_28413030 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[25]));
  AL_DFF_X al_5eade3be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[26]));
  AL_DFF_X al_2ad13761 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[27]));
  AL_DFF_X al_e8fd9177 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[28]));
  AL_DFF_X al_fcbe94a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[29]));
  AL_DFF_X al_81dccbe5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[30]));
  AL_DFF_X al_1d05d28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[31]));
  AL_DFF_X al_fa0a7651 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[32]));
  AL_DFF_X al_1e350978 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[33]));
  AL_DFF_X al_d6c676eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[34]));
  AL_DFF_X al_bb1fbc52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[35]));
  AL_DFF_X al_478abddf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[36]));
  AL_DFF_X al_5d6fa17b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[37]));
  AL_DFF_X al_4a2a548c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[38]));
  AL_DFF_X al_19b33e17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[7]));
  AL_DFF_X al_57ed74a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2ecc3265[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_615b2119[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_2704b644 (
    .a(1'b0),
    .o({al_7581bd0d,open_n167}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_936be3c4 (
    .a(al_7af0d249[8]),
    .b(al_2ecc3265[8]),
    .c(al_7581bd0d),
    .o({al_f01e9810,al_1d982a67[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8d58a6a5 (
    .a(al_7af0d249[9]),
    .b(al_2ecc3265[9]),
    .c(al_f01e9810),
    .o({al_4b0822cb,al_1d982a67[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_30b860f5 (
    .a(al_7af0d249[10]),
    .b(al_2ecc3265[10]),
    .c(al_4b0822cb),
    .o({al_46ca2999,al_1d982a67[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cefe7901 (
    .a(al_7af0d249[11]),
    .b(al_2ecc3265[11]),
    .c(al_46ca2999),
    .o({al_f327e49f,al_1d982a67[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_498ac620 (
    .a(al_7af0d249[12]),
    .b(al_2ecc3265[12]),
    .c(al_f327e49f),
    .o({al_6af99fb0,al_1d982a67[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_823d52c (
    .a(al_7af0d249[13]),
    .b(al_2ecc3265[13]),
    .c(al_6af99fb0),
    .o({al_f9708799,al_1d982a67[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e5c7030d (
    .a(al_7af0d249[14]),
    .b(al_2ecc3265[14]),
    .c(al_f9708799),
    .o({al_ce755696,al_1d982a67[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_253939b9 (
    .a(al_7af0d249[15]),
    .b(al_2ecc3265[15]),
    .c(al_ce755696),
    .o({al_8ceeb1d6,al_1d982a67[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8ca7f1dd (
    .a(al_7af0d249[16]),
    .b(al_2ecc3265[16]),
    .c(al_8ceeb1d6),
    .o({al_56f936a,al_1d982a67[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_126c9a55 (
    .a(al_7af0d249[17]),
    .b(al_2ecc3265[17]),
    .c(al_56f936a),
    .o({al_c17b3665,al_1d982a67[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_961db40 (
    .a(al_7af0d249[18]),
    .b(al_2ecc3265[18]),
    .c(al_c17b3665),
    .o({al_4942e686,al_1d982a67[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_164dbb83 (
    .a(al_7af0d249[19]),
    .b(al_2ecc3265[19]),
    .c(al_4942e686),
    .o({al_fa0cd080,al_1d982a67[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_78f01f82 (
    .a(al_7af0d249[20]),
    .b(al_2ecc3265[20]),
    .c(al_fa0cd080),
    .o({al_b938610a,al_1d982a67[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_51efa356 (
    .a(al_7af0d249[21]),
    .b(al_2ecc3265[21]),
    .c(al_b938610a),
    .o({al_76221ee1,al_1d982a67[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2582d36d (
    .a(al_7af0d249[22]),
    .b(al_2ecc3265[22]),
    .c(al_76221ee1),
    .o({al_73d542b1,al_1d982a67[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_94fbf62f (
    .a(al_7af0d249[23]),
    .b(al_2ecc3265[23]),
    .c(al_73d542b1),
    .o({al_a0e7f496,al_1d982a67[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ae10e38b (
    .a(al_7af0d249[24]),
    .b(al_2ecc3265[24]),
    .c(al_a0e7f496),
    .o({al_5516d10,al_1d982a67[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6db6b6ce (
    .a(al_7af0d249[25]),
    .b(al_2ecc3265[25]),
    .c(al_5516d10),
    .o({al_cade3756,al_1d982a67[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6d962449 (
    .a(al_7af0d249[26]),
    .b(al_2ecc3265[26]),
    .c(al_cade3756),
    .o({al_dc3daad0,al_1d982a67[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_867befa1 (
    .a(al_7af0d249[27]),
    .b(al_2ecc3265[27]),
    .c(al_dc3daad0),
    .o({al_cf98adbf,al_1d982a67[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_af879def (
    .a(al_7af0d249[28]),
    .b(al_2ecc3265[28]),
    .c(al_cf98adbf),
    .o({al_b30ebdf6,al_1d982a67[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_840d4039 (
    .a(al_7af0d249[29]),
    .b(al_2ecc3265[29]),
    .c(al_b30ebdf6),
    .o({al_2258030e,al_1d982a67[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff7a7658 (
    .a(al_7af0d249[30]),
    .b(al_2ecc3265[30]),
    .c(al_2258030e),
    .o({al_8bfba661,al_1d982a67[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d504ad3a (
    .a(al_7af0d249[31]),
    .b(al_2ecc3265[31]),
    .c(al_8bfba661),
    .o({al_9e4c11b8,al_1d982a67[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f3d5ad7b (
    .a(al_7af0d249[32]),
    .b(al_2ecc3265[32]),
    .c(al_9e4c11b8),
    .o({al_7116cd2,al_1d982a67[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_aa96fb8c (
    .a(al_7af0d249[33]),
    .b(al_2ecc3265[33]),
    .c(al_7116cd2),
    .o({al_7c2f83cb,al_1d982a67[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_43daaeef (
    .a(al_7af0d249[34]),
    .b(al_2ecc3265[34]),
    .c(al_7c2f83cb),
    .o({al_689a4219,al_1d982a67[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_45d381f0 (
    .a(al_7af0d249[35]),
    .b(al_2ecc3265[35]),
    .c(al_689a4219),
    .o({al_6d6bb647,al_1d982a67[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ac4a9beb (
    .a(al_7af0d249[36]),
    .b(al_2ecc3265[36]),
    .c(al_6d6bb647),
    .o({al_d9a99e6d,al_1d982a67[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_26ad7161 (
    .a(al_7af0d249[37]),
    .b(al_2ecc3265[37]),
    .c(al_d9a99e6d),
    .o({al_d98a025f,al_1d982a67[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9f7d0af3 (
    .a(al_7af0d249[38]),
    .b(al_2ecc3265[38]),
    .c(al_d98a025f),
    .o({al_6272599f,al_1d982a67[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e5671fee (
    .a(al_7af0d249[39]),
    .b(al_2ecc3265[39]),
    .c(al_6272599f),
    .o({al_c512c49,al_1d982a67[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_18cc1626 (
    .a(al_7af0d249[40]),
    .b(1'b0),
    .c(al_c512c49),
    .o({al_40c30b4d,open_n168}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eca52b4d (
    .a(1'b0),
    .b(1'b1),
    .c(al_40c30b4d),
    .o({open_n169,al_de3e7627}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fb47f7e3 (
    .a(al_7af0d249[10]),
    .b(al_1d982a67[2]),
    .c(al_de3e7627),
    .o(al_d9c08430[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_51b72879 (
    .a(al_7af0d249[11]),
    .b(al_1d982a67[3]),
    .c(al_de3e7627),
    .o(al_d9c08430[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bb41674b (
    .a(al_7af0d249[12]),
    .b(al_1d982a67[4]),
    .c(al_de3e7627),
    .o(al_d9c08430[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_21fa6c6e (
    .a(al_7af0d249[13]),
    .b(al_1d982a67[5]),
    .c(al_de3e7627),
    .o(al_d9c08430[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_18120e3c (
    .a(al_7af0d249[14]),
    .b(al_1d982a67[6]),
    .c(al_de3e7627),
    .o(al_d9c08430[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e62fe763 (
    .a(al_7af0d249[15]),
    .b(al_1d982a67[7]),
    .c(al_de3e7627),
    .o(al_d9c08430[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4a8de6b3 (
    .a(al_7af0d249[16]),
    .b(al_1d982a67[8]),
    .c(al_de3e7627),
    .o(al_d9c08430[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e86c6583 (
    .a(al_7af0d249[17]),
    .b(al_1d982a67[9]),
    .c(al_de3e7627),
    .o(al_d9c08430[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fc1b56f7 (
    .a(al_7af0d249[18]),
    .b(al_1d982a67[10]),
    .c(al_de3e7627),
    .o(al_d9c08430[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_88385740 (
    .a(al_7af0d249[19]),
    .b(al_1d982a67[11]),
    .c(al_de3e7627),
    .o(al_d9c08430[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_31a95722 (
    .a(al_7af0d249[20]),
    .b(al_1d982a67[12]),
    .c(al_de3e7627),
    .o(al_d9c08430[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d31d9d80 (
    .a(al_7af0d249[21]),
    .b(al_1d982a67[13]),
    .c(al_de3e7627),
    .o(al_d9c08430[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c00215d2 (
    .a(al_7af0d249[22]),
    .b(al_1d982a67[14]),
    .c(al_de3e7627),
    .o(al_d9c08430[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bb84d91d (
    .a(al_7af0d249[23]),
    .b(al_1d982a67[15]),
    .c(al_de3e7627),
    .o(al_d9c08430[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_21de10a2 (
    .a(al_7af0d249[24]),
    .b(al_1d982a67[16]),
    .c(al_de3e7627),
    .o(al_d9c08430[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c6393531 (
    .a(al_7af0d249[25]),
    .b(al_1d982a67[17]),
    .c(al_de3e7627),
    .o(al_d9c08430[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1b44f20e (
    .a(al_7af0d249[26]),
    .b(al_1d982a67[18]),
    .c(al_de3e7627),
    .o(al_d9c08430[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_56651036 (
    .a(al_7af0d249[27]),
    .b(al_1d982a67[19]),
    .c(al_de3e7627),
    .o(al_d9c08430[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3d15046 (
    .a(al_7af0d249[28]),
    .b(al_1d982a67[20]),
    .c(al_de3e7627),
    .o(al_d9c08430[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8a2d5974 (
    .a(al_7af0d249[29]),
    .b(al_1d982a67[21]),
    .c(al_de3e7627),
    .o(al_d9c08430[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b995d4ba (
    .a(al_7af0d249[30]),
    .b(al_1d982a67[22]),
    .c(al_de3e7627),
    .o(al_d9c08430[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_531e46c9 (
    .a(al_7af0d249[31]),
    .b(al_1d982a67[23]),
    .c(al_de3e7627),
    .o(al_d9c08430[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bc274ab2 (
    .a(al_7af0d249[32]),
    .b(al_1d982a67[24]),
    .c(al_de3e7627),
    .o(al_d9c08430[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2ffc3487 (
    .a(al_7af0d249[33]),
    .b(al_1d982a67[25]),
    .c(al_de3e7627),
    .o(al_d9c08430[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8b90b901 (
    .a(al_7af0d249[34]),
    .b(al_1d982a67[26]),
    .c(al_de3e7627),
    .o(al_d9c08430[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_aa42d3af (
    .a(al_7af0d249[35]),
    .b(al_1d982a67[27]),
    .c(al_de3e7627),
    .o(al_d9c08430[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_58278aa8 (
    .a(al_7af0d249[36]),
    .b(al_1d982a67[28]),
    .c(al_de3e7627),
    .o(al_d9c08430[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cacc3824 (
    .a(al_7af0d249[37]),
    .b(al_1d982a67[29]),
    .c(al_de3e7627),
    .o(al_d9c08430[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c08e6570 (
    .a(al_7af0d249[38]),
    .b(al_1d982a67[30]),
    .c(al_de3e7627),
    .o(al_d9c08430[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_71546d65 (
    .a(al_7af0d249[39]),
    .b(al_1d982a67[31]),
    .c(al_de3e7627),
    .o(al_d9c08430[39]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_56ca5c23 (
    .a(al_7af0d249[8]),
    .b(al_1d982a67[0]),
    .c(al_de3e7627),
    .o(al_d9c08430[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9a3ae1b8 (
    .a(al_7af0d249[9]),
    .b(al_1d982a67[1]),
    .c(al_de3e7627),
    .o(al_d9c08430[9]));
  AL_DFF_X al_d231dfce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7af0d249[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[0]));
  AL_DFF_X al_c887eba4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[9]));
  AL_DFF_X al_6588317f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[10]));
  AL_DFF_X al_3560567f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[11]));
  AL_DFF_X al_55926c03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[12]));
  AL_DFF_X al_d410f217 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[13]));
  AL_DFF_X al_83ec1453 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[14]));
  AL_DFF_X al_e4629127 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[15]));
  AL_DFF_X al_26e879bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[16]));
  AL_DFF_X al_55a9183d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[17]));
  AL_DFF_X al_70432270 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[18]));
  AL_DFF_X al_3c5c3bf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7af0d249[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[1]));
  AL_DFF_X al_ab543f44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[19]));
  AL_DFF_X al_ecdc60df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[20]));
  AL_DFF_X al_65792b32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[21]));
  AL_DFF_X al_6bff2632 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[22]));
  AL_DFF_X al_e17908c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[23]));
  AL_DFF_X al_bc564939 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[24]));
  AL_DFF_X al_c930a2e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[25]));
  AL_DFF_X al_1d4c4f47 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[26]));
  AL_DFF_X al_1020e795 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[27]));
  AL_DFF_X al_22db711c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[28]));
  AL_DFF_X al_faf12c7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7af0d249[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[2]));
  AL_DFF_X al_dce2c5ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[29]));
  AL_DFF_X al_c3fd716d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[30]));
  AL_DFF_X al_3044694a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[31]));
  AL_DFF_X al_c0f165f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[32]));
  AL_DFF_X al_649b3c8f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[33]));
  AL_DFF_X al_243f09e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[34]));
  AL_DFF_X al_bf8799f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[35]));
  AL_DFF_X al_d50abc6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[36]));
  AL_DFF_X al_9a72c743 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[37]));
  AL_DFF_X al_aa4da4f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[38]));
  AL_DFF_X al_80f1f5a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7af0d249[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[3]));
  AL_DFF_X al_a853ef6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[39]));
  AL_DFF_X al_d6c510ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7af0d249[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[4]));
  AL_DFF_X al_2d6cb65c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7af0d249[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[5]));
  AL_DFF_X al_9bcf9550 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7af0d249[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[6]));
  AL_DFF_X al_811f2d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7af0d249[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[7]));
  AL_DFF_X al_990bacfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d9c08430[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ce3b275[8]));
  AL_DFF_X al_314a9cd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_de3e7627),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[0]));
  AL_DFF_X al_1ea8ad71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[9]));
  AL_DFF_X al_ed5e87f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[10]));
  AL_DFF_X al_463c1455 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[11]));
  AL_DFF_X al_f90f36eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[12]));
  AL_DFF_X al_e5c5f2f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[13]));
  AL_DFF_X al_547b7e63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[14]));
  AL_DFF_X al_c58c4aea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[15]));
  AL_DFF_X al_86a31641 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[16]));
  AL_DFF_X al_91e3373e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[17]));
  AL_DFF_X al_3451a7bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[18]));
  AL_DFF_X al_f48ff60c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[1]));
  AL_DFF_X al_b8cb84af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[19]));
  AL_DFF_X al_5ba24f5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[20]));
  AL_DFF_X al_20f24576 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[21]));
  AL_DFF_X al_be44438e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[22]));
  AL_DFF_X al_a6d76b2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[23]));
  AL_DFF_X al_c818df74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[24]));
  AL_DFF_X al_8ad45735 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[25]));
  AL_DFF_X al_3cd09252 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[26]));
  AL_DFF_X al_e2f6f95a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[27]));
  AL_DFF_X al_8ef89d11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[28]));
  AL_DFF_X al_3be16670 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[2]));
  AL_DFF_X al_6b52a3ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[29]));
  AL_DFF_X al_4aa66622 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[30]));
  AL_DFF_X al_1cc50bee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[31]));
  AL_DFF_X al_19c9b251 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[32]));
  AL_DFF_X al_7870e5f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[33]));
  AL_DFF_X al_1f557b52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[34]));
  AL_DFF_X al_e9780f00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[35]));
  AL_DFF_X al_9312c378 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[36]));
  AL_DFF_X al_9493b03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[37]));
  AL_DFF_X al_e91177b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[38]));
  AL_DFF_X al_9a0747d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[3]));
  AL_DFF_X al_1a1ebc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[39]));
  AL_DFF_X al_31aa1bfe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[4]));
  AL_DFF_X al_dded1598 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[5]));
  AL_DFF_X al_ba93379d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[6]));
  AL_DFF_X al_df0c3fa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[7]));
  AL_DFF_X al_e7787cdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b6775e93[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_56efbba9[8]));
  AL_DFF_X al_d3b07a22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44882eca[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f336c405[0]));
  AL_DFF_X al_b79d8302 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[43]));
  AL_DFF_X al_3b200631 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[44]));
  AL_DFF_X al_995d2c96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[45]));
  AL_DFF_X al_d2e46076 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[46]));
  AL_DFF_X al_5895eba4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[47]));
  AL_DFF_X al_761ee1f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[48]));
  AL_DFF_X al_ed810f78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[49]));
  AL_DFF_X al_4b59d924 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[50]));
  AL_DFF_X al_46960228 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[51]));
  AL_DFF_X al_a34ec6e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[52]));
  AL_DFF_X al_ea2dac2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[53]));
  AL_DFF_X al_30b87125 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[54]));
  AL_DFF_X al_2abf5269 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[55]));
  AL_DFF_X al_1d810297 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[56]));
  AL_DFF_X al_37ca961a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[57]));
  AL_DFF_X al_b8d7a90c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[58]));
  AL_DFF_X al_e2c17710 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[59]));
  AL_DFF_X al_20ef2f11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[60]));
  AL_DFF_X al_ce90d7c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[61]));
  AL_DFF_X al_24c6e74f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[62]));
  AL_DFF_X al_d53beca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[63]));
  AL_DFF_X al_9d8c6bfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[64]));
  AL_DFF_X al_709d6b8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[65]));
  AL_DFF_X al_23533eb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[66]));
  AL_DFF_X al_b27220a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[67]));
  AL_DFF_X al_d858d7db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[68]));
  AL_DFF_X al_ddee2f21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[69]));
  AL_DFF_X al_83f53d26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[70]));
  AL_DFF_X al_dd9f120b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[71]));
  AL_DFF_X al_a643c27e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[72]));
  AL_DFF_X al_d842fbc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[73]));
  AL_DFF_X al_dadd0006 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b052c226[75]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_28202fa7[74]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    al_3b7b1f10 (
    .a(al_7d13d94f),
    .b(al_626a930b),
    .c(al_ab96385b),
    .o(al_b2787015));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((~D*A))*~(E)*~(F)+~(B)*~(C)*~((~D*A))*E*~(F)+B*~(C)*~((~D*A))*E*~(F)+~(B)*~(C)*(~D*A)*E*~(F)+~(B)*~(C)*~((~D*A))*~(E)*F+B*~(C)*~((~D*A))*~(E)*F+~(B)*C*~((~D*A))*~(E)*F+~(B)*~(C)*(~D*A)*~(E)*F+B*~(C)*(~D*A)*~(E)*F+~(B)*~(C)*~((~D*A))*E*F+B*~(C)*~((~D*A))*E*F+~(B)*C*~((~D*A))*E*F+B*C*~((~D*A))*E*F+~(B)*~(C)*(~D*A)*E*F+B*~(C)*(~D*A)*E*F+~(B)*C*(~D*A)*E*F)"),
    .INIT(64'hff7f3f1f0f070301))
    al_1aecd3bc (
    .a(al_b052c226[44]),
    .b(al_b052c226[45]),
    .c(al_b052c226[46]),
    .d(al_592f1b09[44]),
    .e(al_592f1b09[45]),
    .f(al_592f1b09[46]),
    .o(al_92ccaa05));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_5a6fe739 (
    .a(al_b052c226[61]),
    .b(al_b052c226[62]),
    .c(al_b052c226[65]),
    .d(al_b052c226[66]),
    .e(al_b052c226[68]),
    .f(al_b052c226[71]),
    .o(al_3bcfaff1));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_2e66739 (
    .a(al_b052c226[49]),
    .b(al_b052c226[50]),
    .c(al_b052c226[52]),
    .d(al_b052c226[55]),
    .e(al_b052c226[56]),
    .f(al_b052c226[59]),
    .o(al_4059e403));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    al_b0fb52ad (
    .a(al_3bcfaff1),
    .b(al_4059e403),
    .o(al_ab96385b));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*C*B*~A))"),
    .INIT(32'hbfff4000))
    al_a2a70cd0 (
    .a(al_7d13d94f),
    .b(al_626a930b),
    .c(al_ab96385b),
    .d(al_b052c226[44]),
    .e(al_592f1b09[44]),
    .o(al_8c015879[44]));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*B*C)"),
    .INIT(8'h4d))
    al_9c9b16b4 (
    .a(al_92ccaa05),
    .b(al_b052c226[47]),
    .c(al_592f1b09[47]),
    .o(al_7d13d94f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_6ff36723 (
    .a(al_b052c226[69]),
    .b(al_b052c226[70]),
    .c(al_b052c226[72]),
    .d(al_b052c226[73]),
    .e(al_b052c226[74]),
    .f(al_b052c226[75]),
    .o(al_b458e911));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_b5180229 (
    .a(al_b052c226[57]),
    .b(al_b052c226[58]),
    .c(al_b052c226[60]),
    .d(al_b052c226[63]),
    .e(al_b052c226[64]),
    .f(al_b052c226[67]),
    .o(al_f5397afe));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*B*A)"),
    .INIT(64'h0000000000000008))
    al_55b2bb57 (
    .a(al_b458e911),
    .b(al_f5397afe),
    .c(al_b052c226[48]),
    .d(al_b052c226[51]),
    .e(al_b052c226[53]),
    .f(al_b052c226[54]),
    .o(al_626a930b));
  AL_MAP_LUT5 #(
    .EQN("(B*A*(D@(~E*C)))"),
    .INIT(32'h88000880))
    al_1093a0e2 (
    .a(al_3bcfaff1),
    .b(al_4059e403),
    .c(al_b052c226[44]),
    .d(al_b052c226[45]),
    .e(al_592f1b09[44]),
    .o(al_12b84efd));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*B*~A))"),
    .INIT(16'hbf40))
    al_f248a313 (
    .a(al_7d13d94f),
    .b(al_626a930b),
    .c(al_12b84efd),
    .d(al_592f1b09[45]),
    .o(al_8c015879[45]));
  AL_MAP_LUT5 #(
    .EQN("(C@(B*~((~D*A))*~(E)+~(B)*(~D*A)*~(E)+B*(~D*A)*~(E)+B*(~D*A)*E))"),
    .INIT(32'hf0783c1e))
    al_4e8e7c8f (
    .a(al_b052c226[44]),
    .b(al_b052c226[45]),
    .c(al_b052c226[46]),
    .d(al_592f1b09[44]),
    .e(al_592f1b09[45]),
    .o(al_40670ee4));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*C*B*~A))"),
    .INIT(32'hbfff4000))
    al_4f9326e8 (
    .a(al_7d13d94f),
    .b(al_626a930b),
    .c(al_ab96385b),
    .d(al_40670ee4),
    .e(al_592f1b09[46]),
    .o(al_8c015879[46]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(B*A*~(D@C)))"),
    .INIT(32'h7ff70000))
    al_fcb4ba27 (
    .a(al_626a930b),
    .b(al_ab96385b),
    .c(al_92ccaa05),
    .d(al_b052c226[47]),
    .e(al_592f1b09[47]),
    .o(al_8c015879[47]));
  AL_DFF_X al_86e9db3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[0]));
  AL_DFF_X al_9781634b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[9]));
  AL_DFF_X al_6b03f0d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[10]));
  AL_DFF_X al_9bb317a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[11]));
  AL_DFF_X al_fb93ead8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[12]));
  AL_DFF_X al_64415bdb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[13]));
  AL_DFF_X al_c27ef722 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[14]));
  AL_DFF_X al_152877f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[15]));
  AL_DFF_X al_b5afc7e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[16]));
  AL_DFF_X al_30ab2183 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[17]));
  AL_DFF_X al_cba85855 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[18]));
  AL_DFF_X al_36402053 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[1]));
  AL_DFF_X al_2b7dfadf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[19]));
  AL_DFF_X al_8d1cee72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[20]));
  AL_DFF_X al_8c32f1c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[21]));
  AL_DFF_X al_38a7a2f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[22]));
  AL_DFF_X al_ea342da5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[23]));
  AL_DFF_X al_25967989 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[24]));
  AL_DFF_X al_307b0033 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[25]));
  AL_DFF_X al_b63216b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[26]));
  AL_DFF_X al_a899fcbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[27]));
  AL_DFF_X al_21320ba3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[28]));
  AL_DFF_X al_113f7fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[2]));
  AL_DFF_X al_3634fc15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[29]));
  AL_DFF_X al_69b783ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[30]));
  AL_DFF_X al_e1d51dca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[31]));
  AL_DFF_X al_4491657f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[32]));
  AL_DFF_X al_39070cdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[33]));
  AL_DFF_X al_f876df13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[34]));
  AL_DFF_X al_cc9cec3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[35]));
  AL_DFF_X al_ebad2beb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[36]));
  AL_DFF_X al_a6bc2c04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[37]));
  AL_DFF_X al_51e4ee4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[38]));
  AL_DFF_X al_ac3cf438 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[3]));
  AL_DFF_X al_62980d6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[39]));
  AL_DFF_X al_c832177f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[40]));
  AL_DFF_X al_dcec40bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[41]));
  AL_DFF_X al_c44ae4c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[42]));
  AL_DFF_X al_2cbf3751 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[43]));
  AL_DFF_X al_75130f02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c015879[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[44]));
  AL_DFF_X al_7102ad96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c015879[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[45]));
  AL_DFF_X al_62a12f1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c015879[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[46]));
  AL_DFF_X al_64448bba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8c015879[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[47]));
  AL_DFF_X al_121d90f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[4]));
  AL_DFF_X al_bd4611bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[5]));
  AL_DFF_X al_bc8790b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[6]));
  AL_DFF_X al_644842b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[7]));
  AL_DFF_X al_32d7571 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_592f1b09[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1d4399b1[8]));
  AL_DFF_X al_4ad54e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b2787015),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_917df14b[0]));
  AL_DFF_X al_f307e68b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b18b7cbb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_917df14b[1]));
  AL_DFF_X al_11748906 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b18b7cbb[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_917df14b[2]));
  AL_DFF_X al_1f4fa5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b18b7cbb[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_917df14b[3]));
  AL_DFF_X al_3ff12f07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5bcbf559[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_16eefd24[0]));
  AL_DFF_X al_693c0f87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[9]));
  AL_DFF_X al_8eda5251 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[10]));
  AL_DFF_X al_fe9b0f0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[11]));
  AL_DFF_X al_312fcdd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[12]));
  AL_DFF_X al_9deab9cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[13]));
  AL_DFF_X al_a9d604e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[14]));
  AL_DFF_X al_ab5d0b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[15]));
  AL_DFF_X al_be8d0355 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[16]));
  AL_DFF_X al_f38bc011 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[17]));
  AL_DFF_X al_2eb315b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[18]));
  AL_DFF_X al_b24ddd6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[19]));
  AL_DFF_X al_4b1328d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[20]));
  AL_DFF_X al_32b32e14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[21]));
  AL_DFF_X al_4d394b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[22]));
  AL_DFF_X al_f4723a80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[23]));
  AL_DFF_X al_dd97123e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[24]));
  AL_DFF_X al_c43921ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[25]));
  AL_DFF_X al_6ec41f5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[26]));
  AL_DFF_X al_3c457c2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[27]));
  AL_DFF_X al_1a33428 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[28]));
  AL_DFF_X al_b4067bc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[29]));
  AL_DFF_X al_c7c58acf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[30]));
  AL_DFF_X al_39c613a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[31]));
  AL_DFF_X al_8f9b1864 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[32]));
  AL_DFF_X al_d6fb0960 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[33]));
  AL_DFF_X al_eb9aa2d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[34]));
  AL_DFF_X al_891030a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[35]));
  AL_DFF_X al_d9b12eec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[36]));
  AL_DFF_X al_68ba2fa4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[37]));
  AL_DFF_X al_2ac74e2e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[6]));
  AL_DFF_X al_29053179 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[7]));
  AL_DFF_X al_bb21e43f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_615b2119[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_aa3e519e[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_85a4bc22 (
    .a(1'b0),
    .o({al_e23a271f,open_n172}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a7e6059 (
    .a(al_ce3b275[7]),
    .b(al_615b2119[7]),
    .c(al_e23a271f),
    .o({al_eed33fc3,al_79977513[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fd023b0d (
    .a(al_ce3b275[8]),
    .b(al_615b2119[8]),
    .c(al_eed33fc3),
    .o({al_7e086938,al_79977513[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b6f42af (
    .a(al_ce3b275[9]),
    .b(al_615b2119[9]),
    .c(al_7e086938),
    .o({al_4ebf21a,al_79977513[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8aa388a7 (
    .a(al_ce3b275[10]),
    .b(al_615b2119[10]),
    .c(al_4ebf21a),
    .o({al_f74ec05f,al_79977513[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_947b917 (
    .a(al_ce3b275[11]),
    .b(al_615b2119[11]),
    .c(al_f74ec05f),
    .o({al_b1a4aa4,al_79977513[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cac68a51 (
    .a(al_ce3b275[12]),
    .b(al_615b2119[12]),
    .c(al_b1a4aa4),
    .o({al_98dec4e,al_79977513[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_99660cc2 (
    .a(al_ce3b275[13]),
    .b(al_615b2119[13]),
    .c(al_98dec4e),
    .o({al_2825c36a,al_79977513[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b05f5683 (
    .a(al_ce3b275[14]),
    .b(al_615b2119[14]),
    .c(al_2825c36a),
    .o({al_ca256ef5,al_79977513[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4b9d1fc7 (
    .a(al_ce3b275[15]),
    .b(al_615b2119[15]),
    .c(al_ca256ef5),
    .o({al_cac22815,al_79977513[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8c5a91b7 (
    .a(al_ce3b275[16]),
    .b(al_615b2119[16]),
    .c(al_cac22815),
    .o({al_7b366c25,al_79977513[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c3764128 (
    .a(al_ce3b275[17]),
    .b(al_615b2119[17]),
    .c(al_7b366c25),
    .o({al_306af3cf,al_79977513[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67604e75 (
    .a(al_ce3b275[18]),
    .b(al_615b2119[18]),
    .c(al_306af3cf),
    .o({al_4957c6a5,al_79977513[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c7eb7372 (
    .a(al_ce3b275[19]),
    .b(al_615b2119[19]),
    .c(al_4957c6a5),
    .o({al_8a47c612,al_79977513[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_19d5b1ef (
    .a(al_ce3b275[20]),
    .b(al_615b2119[20]),
    .c(al_8a47c612),
    .o({al_f65c10,al_79977513[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_42b19f46 (
    .a(al_ce3b275[21]),
    .b(al_615b2119[21]),
    .c(al_f65c10),
    .o({al_6a66d91e,al_79977513[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2ace5dda (
    .a(al_ce3b275[22]),
    .b(al_615b2119[22]),
    .c(al_6a66d91e),
    .o({al_bcbd4e1b,al_79977513[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68b10a87 (
    .a(al_ce3b275[23]),
    .b(al_615b2119[23]),
    .c(al_bcbd4e1b),
    .o({al_792f9fb1,al_79977513[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_baaa4a68 (
    .a(al_ce3b275[24]),
    .b(al_615b2119[24]),
    .c(al_792f9fb1),
    .o({al_1f9c650e,al_79977513[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e99a601f (
    .a(al_ce3b275[25]),
    .b(al_615b2119[25]),
    .c(al_1f9c650e),
    .o({al_e88204f,al_79977513[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5f0dda22 (
    .a(al_ce3b275[26]),
    .b(al_615b2119[26]),
    .c(al_e88204f),
    .o({al_c435b5e6,al_79977513[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a5efa223 (
    .a(al_ce3b275[27]),
    .b(al_615b2119[27]),
    .c(al_c435b5e6),
    .o({al_13c84cc8,al_79977513[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6a730672 (
    .a(al_ce3b275[28]),
    .b(al_615b2119[28]),
    .c(al_13c84cc8),
    .o({al_21c2c54f,al_79977513[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e7f2bc7d (
    .a(al_ce3b275[29]),
    .b(al_615b2119[29]),
    .c(al_21c2c54f),
    .o({al_fe48089b,al_79977513[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5aa57ad7 (
    .a(al_ce3b275[30]),
    .b(al_615b2119[30]),
    .c(al_fe48089b),
    .o({al_fe0b2c2e,al_79977513[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7a9e140a (
    .a(al_ce3b275[31]),
    .b(al_615b2119[31]),
    .c(al_fe0b2c2e),
    .o({al_8b619c3b,al_79977513[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4f058c6d (
    .a(al_ce3b275[32]),
    .b(al_615b2119[32]),
    .c(al_8b619c3b),
    .o({al_a522c3d4,al_79977513[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_774ebe73 (
    .a(al_ce3b275[33]),
    .b(al_615b2119[33]),
    .c(al_a522c3d4),
    .o({al_e347376a,al_79977513[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a6b0d1a9 (
    .a(al_ce3b275[34]),
    .b(al_615b2119[34]),
    .c(al_e347376a),
    .o({al_28f6cbc1,al_79977513[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_544deb8a (
    .a(al_ce3b275[35]),
    .b(al_615b2119[35]),
    .c(al_28f6cbc1),
    .o({al_17617f0f,al_79977513[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_97826cc9 (
    .a(al_ce3b275[36]),
    .b(al_615b2119[36]),
    .c(al_17617f0f),
    .o({al_510c2901,al_79977513[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_14ddc944 (
    .a(al_ce3b275[37]),
    .b(al_615b2119[37]),
    .c(al_510c2901),
    .o({al_8aca8bdd,al_79977513[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9bcab770 (
    .a(al_ce3b275[38]),
    .b(al_615b2119[38]),
    .c(al_8aca8bdd),
    .o({al_94c5d51b,al_79977513[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_32d8a393 (
    .a(al_ce3b275[39]),
    .b(1'b0),
    .c(al_94c5d51b),
    .o({al_ec8c91da,open_n173}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_53748320 (
    .a(1'b0),
    .b(1'b1),
    .c(al_ec8c91da),
    .o({open_n174,al_a1bb6a32}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6bafebba (
    .a(al_ce3b275[10]),
    .b(al_79977513[3]),
    .c(al_a1bb6a32),
    .o(al_92415709[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ed680f64 (
    .a(al_ce3b275[11]),
    .b(al_79977513[4]),
    .c(al_a1bb6a32),
    .o(al_92415709[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_836c9272 (
    .a(al_ce3b275[12]),
    .b(al_79977513[5]),
    .c(al_a1bb6a32),
    .o(al_92415709[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b40fbca7 (
    .a(al_ce3b275[13]),
    .b(al_79977513[6]),
    .c(al_a1bb6a32),
    .o(al_92415709[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fd33a3b0 (
    .a(al_ce3b275[14]),
    .b(al_79977513[7]),
    .c(al_a1bb6a32),
    .o(al_92415709[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_af26f540 (
    .a(al_ce3b275[15]),
    .b(al_79977513[8]),
    .c(al_a1bb6a32),
    .o(al_92415709[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5fea570 (
    .a(al_ce3b275[16]),
    .b(al_79977513[9]),
    .c(al_a1bb6a32),
    .o(al_92415709[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_45916ff5 (
    .a(al_ce3b275[17]),
    .b(al_79977513[10]),
    .c(al_a1bb6a32),
    .o(al_92415709[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_10fdb491 (
    .a(al_ce3b275[18]),
    .b(al_79977513[11]),
    .c(al_a1bb6a32),
    .o(al_92415709[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d5e6e4c9 (
    .a(al_ce3b275[19]),
    .b(al_79977513[12]),
    .c(al_a1bb6a32),
    .o(al_92415709[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c9536a94 (
    .a(al_ce3b275[20]),
    .b(al_79977513[13]),
    .c(al_a1bb6a32),
    .o(al_92415709[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_be5f6f58 (
    .a(al_ce3b275[21]),
    .b(al_79977513[14]),
    .c(al_a1bb6a32),
    .o(al_92415709[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_740eb3cc (
    .a(al_ce3b275[22]),
    .b(al_79977513[15]),
    .c(al_a1bb6a32),
    .o(al_92415709[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d2e2b00 (
    .a(al_ce3b275[23]),
    .b(al_79977513[16]),
    .c(al_a1bb6a32),
    .o(al_92415709[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_49f11be6 (
    .a(al_ce3b275[24]),
    .b(al_79977513[17]),
    .c(al_a1bb6a32),
    .o(al_92415709[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4dc96c5f (
    .a(al_ce3b275[25]),
    .b(al_79977513[18]),
    .c(al_a1bb6a32),
    .o(al_92415709[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_59cf2081 (
    .a(al_ce3b275[26]),
    .b(al_79977513[19]),
    .c(al_a1bb6a32),
    .o(al_92415709[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_669327c3 (
    .a(al_ce3b275[27]),
    .b(al_79977513[20]),
    .c(al_a1bb6a32),
    .o(al_92415709[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8f644ee1 (
    .a(al_ce3b275[28]),
    .b(al_79977513[21]),
    .c(al_a1bb6a32),
    .o(al_92415709[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_44a1f566 (
    .a(al_ce3b275[29]),
    .b(al_79977513[22]),
    .c(al_a1bb6a32),
    .o(al_92415709[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e5bed236 (
    .a(al_ce3b275[30]),
    .b(al_79977513[23]),
    .c(al_a1bb6a32),
    .o(al_92415709[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_93910ff8 (
    .a(al_ce3b275[31]),
    .b(al_79977513[24]),
    .c(al_a1bb6a32),
    .o(al_92415709[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b00d3cf2 (
    .a(al_ce3b275[32]),
    .b(al_79977513[25]),
    .c(al_a1bb6a32),
    .o(al_92415709[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_69de3d12 (
    .a(al_ce3b275[33]),
    .b(al_79977513[26]),
    .c(al_a1bb6a32),
    .o(al_92415709[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e14a37db (
    .a(al_ce3b275[34]),
    .b(al_79977513[27]),
    .c(al_a1bb6a32),
    .o(al_92415709[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ebf477f4 (
    .a(al_ce3b275[35]),
    .b(al_79977513[28]),
    .c(al_a1bb6a32),
    .o(al_92415709[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e2778e22 (
    .a(al_ce3b275[36]),
    .b(al_79977513[29]),
    .c(al_a1bb6a32),
    .o(al_92415709[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ab0584bd (
    .a(al_ce3b275[37]),
    .b(al_79977513[30]),
    .c(al_a1bb6a32),
    .o(al_92415709[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c051d9dc (
    .a(al_ce3b275[38]),
    .b(al_79977513[31]),
    .c(al_a1bb6a32),
    .o(al_92415709[38]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9a3b1a20 (
    .a(al_ce3b275[7]),
    .b(al_79977513[0]),
    .c(al_a1bb6a32),
    .o(al_92415709[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_49cb43eb (
    .a(al_ce3b275[8]),
    .b(al_79977513[1]),
    .c(al_a1bb6a32),
    .o(al_92415709[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5cd7fec2 (
    .a(al_ce3b275[9]),
    .b(al_79977513[2]),
    .c(al_a1bb6a32),
    .o(al_92415709[9]));
  AL_DFF_X al_22de739 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce3b275[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[0]));
  AL_DFF_X al_c69c8e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[9]));
  AL_DFF_X al_b96719ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[10]));
  AL_DFF_X al_b0795a10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[11]));
  AL_DFF_X al_730ca21e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[12]));
  AL_DFF_X al_f0891dd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[13]));
  AL_DFF_X al_92da3b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[14]));
  AL_DFF_X al_55a174ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[15]));
  AL_DFF_X al_cf617560 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[16]));
  AL_DFF_X al_1686e8e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[17]));
  AL_DFF_X al_9b771d55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[18]));
  AL_DFF_X al_c7cef16e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce3b275[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[1]));
  AL_DFF_X al_210ec171 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[19]));
  AL_DFF_X al_fe78fbc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[20]));
  AL_DFF_X al_a7977a79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[21]));
  AL_DFF_X al_ccb400c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[22]));
  AL_DFF_X al_2730cdb0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[23]));
  AL_DFF_X al_6ec787be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[24]));
  AL_DFF_X al_8cf071ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[25]));
  AL_DFF_X al_21d4625c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[26]));
  AL_DFF_X al_3c2e02fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[27]));
  AL_DFF_X al_7504e264 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[28]));
  AL_DFF_X al_30009153 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce3b275[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[2]));
  AL_DFF_X al_c2b55a27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[29]));
  AL_DFF_X al_a0451767 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[30]));
  AL_DFF_X al_545e214b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[31]));
  AL_DFF_X al_4391203b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[32]));
  AL_DFF_X al_5fe51d76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[33]));
  AL_DFF_X al_46f87198 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[34]));
  AL_DFF_X al_9d8bcb64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[35]));
  AL_DFF_X al_53dfa7bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[36]));
  AL_DFF_X al_644a14b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[37]));
  AL_DFF_X al_f591c37e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[38]));
  AL_DFF_X al_bfce5c63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce3b275[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[3]));
  AL_DFF_X al_540a311f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce3b275[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[4]));
  AL_DFF_X al_ca5e3c5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce3b275[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[5]));
  AL_DFF_X al_46641fd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce3b275[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[6]));
  AL_DFF_X al_58517639 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[7]));
  AL_DFF_X al_df23030a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_92415709[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f8daefdd[8]));
  AL_DFF_X al_e925eb5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_a1bb6a32),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[0]));
  AL_DFF_X al_bdb7d525 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[9]));
  AL_DFF_X al_9c58e579 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[10]));
  AL_DFF_X al_eee7353c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[11]));
  AL_DFF_X al_ff748c77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[12]));
  AL_DFF_X al_ce9e8fbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[13]));
  AL_DFF_X al_3ce1618e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[14]));
  AL_DFF_X al_8b8d611a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[15]));
  AL_DFF_X al_5de729cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[16]));
  AL_DFF_X al_842ec08d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[17]));
  AL_DFF_X al_724e7b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[18]));
  AL_DFF_X al_991db7dd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[1]));
  AL_DFF_X al_e5139954 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[19]));
  AL_DFF_X al_960192a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[20]));
  AL_DFF_X al_a795c268 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[21]));
  AL_DFF_X al_58a2cef1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[22]));
  AL_DFF_X al_a3602b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[23]));
  AL_DFF_X al_a5c1815d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[24]));
  AL_DFF_X al_c4eda67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[25]));
  AL_DFF_X al_d536c1ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[26]));
  AL_DFF_X al_f4baf849 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[27]));
  AL_DFF_X al_5b4059ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[28]));
  AL_DFF_X al_edded638 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[2]));
  AL_DFF_X al_d7fa9615 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[29]));
  AL_DFF_X al_efc23e00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[30]));
  AL_DFF_X al_bdc76a7a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[31]));
  AL_DFF_X al_b2d55898 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[32]));
  AL_DFF_X al_4148a085 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[33]));
  AL_DFF_X al_d91f64e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[34]));
  AL_DFF_X al_2cc0c290 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[35]));
  AL_DFF_X al_fb747d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[36]));
  AL_DFF_X al_7a7eb955 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[37]));
  AL_DFF_X al_b7772511 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[38]));
  AL_DFF_X al_35876ebf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[3]));
  AL_DFF_X al_d5122abc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[39]));
  AL_DFF_X al_ae846c45 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[40]));
  AL_DFF_X al_af316b1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[4]));
  AL_DFF_X al_147cae2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[5]));
  AL_DFF_X al_abf82517 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[6]));
  AL_DFF_X al_b22ab5d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[7]));
  AL_DFF_X al_10294f51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_56efbba9[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3357c8f6[8]));
  AL_DFF_X al_99b1d1c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_16eefd24[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_993138f9[0]));
  AL_DFF_X al_fc7b19f3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[9]));
  AL_DFF_X al_afb409fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[10]));
  AL_DFF_X al_d5ed275a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[11]));
  AL_DFF_X al_d1eeaea9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[12]));
  AL_DFF_X al_d61e7254 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[13]));
  AL_DFF_X al_789042c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[14]));
  AL_DFF_X al_5bd522ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[15]));
  AL_DFF_X al_15621d7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[16]));
  AL_DFF_X al_2a0533c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[17]));
  AL_DFF_X al_24c48c2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[18]));
  AL_DFF_X al_7f72f72f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[19]));
  AL_DFF_X al_4612ce33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[20]));
  AL_DFF_X al_537531ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[21]));
  AL_DFF_X al_52c8f3fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[22]));
  AL_DFF_X al_61f18d0a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[23]));
  AL_DFF_X al_d6c05ffa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[24]));
  AL_DFF_X al_94154e71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[25]));
  AL_DFF_X al_7df9f6bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[26]));
  AL_DFF_X al_9c3617ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[27]));
  AL_DFF_X al_11ecdc54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[28]));
  AL_DFF_X al_134b02ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[29]));
  AL_DFF_X al_acaf2b9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[30]));
  AL_DFF_X al_fcfb01d1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[31]));
  AL_DFF_X al_6d48bf7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[32]));
  AL_DFF_X al_c0a7a093 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[33]));
  AL_DFF_X al_cdcf5586 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[34]));
  AL_DFF_X al_3e6a8cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[35]));
  AL_DFF_X al_c2049239 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[36]));
  AL_DFF_X al_1d2eb9fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[5]));
  AL_DFF_X al_f1b02e3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[6]));
  AL_DFF_X al_d656a0f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[7]));
  AL_DFF_X al_611db5b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_aa3e519e[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5e4a13f0[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_e66df217 (
    .a(1'b0),
    .o({al_ac09860,open_n177}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_921dafaa (
    .a(al_f8daefdd[6]),
    .b(al_aa3e519e[6]),
    .c(al_ac09860),
    .o({al_8818311f,al_a972f2b7[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fbd22be3 (
    .a(al_f8daefdd[7]),
    .b(al_aa3e519e[7]),
    .c(al_8818311f),
    .o({al_189a7687,al_a972f2b7[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bb5917e7 (
    .a(al_f8daefdd[8]),
    .b(al_aa3e519e[8]),
    .c(al_189a7687),
    .o({al_b94ff95a,al_a972f2b7[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ca8f8b60 (
    .a(al_f8daefdd[9]),
    .b(al_aa3e519e[9]),
    .c(al_b94ff95a),
    .o({al_1a56b969,al_a972f2b7[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d65199a6 (
    .a(al_f8daefdd[10]),
    .b(al_aa3e519e[10]),
    .c(al_1a56b969),
    .o({al_5971bdb0,al_a972f2b7[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_724d0102 (
    .a(al_f8daefdd[11]),
    .b(al_aa3e519e[11]),
    .c(al_5971bdb0),
    .o({al_a1353883,al_a972f2b7[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_65e7e39c (
    .a(al_f8daefdd[12]),
    .b(al_aa3e519e[12]),
    .c(al_a1353883),
    .o({al_a8675d43,al_a972f2b7[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2969412b (
    .a(al_f8daefdd[13]),
    .b(al_aa3e519e[13]),
    .c(al_a8675d43),
    .o({al_2dcd8322,al_a972f2b7[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1e2cf43b (
    .a(al_f8daefdd[14]),
    .b(al_aa3e519e[14]),
    .c(al_2dcd8322),
    .o({al_1e9d53ff,al_a972f2b7[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ec95dc26 (
    .a(al_f8daefdd[15]),
    .b(al_aa3e519e[15]),
    .c(al_1e9d53ff),
    .o({al_a3e2ac47,al_a972f2b7[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_947babf4 (
    .a(al_f8daefdd[16]),
    .b(al_aa3e519e[16]),
    .c(al_a3e2ac47),
    .o({al_da3e5716,al_a972f2b7[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_af058393 (
    .a(al_f8daefdd[17]),
    .b(al_aa3e519e[17]),
    .c(al_da3e5716),
    .o({al_6b874685,al_a972f2b7[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cff83812 (
    .a(al_f8daefdd[18]),
    .b(al_aa3e519e[18]),
    .c(al_6b874685),
    .o({al_ab74a1e3,al_a972f2b7[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bba1b04b (
    .a(al_f8daefdd[19]),
    .b(al_aa3e519e[19]),
    .c(al_ab74a1e3),
    .o({al_6c10ec91,al_a972f2b7[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bd8525e2 (
    .a(al_f8daefdd[20]),
    .b(al_aa3e519e[20]),
    .c(al_6c10ec91),
    .o({al_c829298,al_a972f2b7[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c55213ff (
    .a(al_f8daefdd[21]),
    .b(al_aa3e519e[21]),
    .c(al_c829298),
    .o({al_88013228,al_a972f2b7[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6d79dcd8 (
    .a(al_f8daefdd[22]),
    .b(al_aa3e519e[22]),
    .c(al_88013228),
    .o({al_ebe24e3d,al_a972f2b7[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_23164bfc (
    .a(al_f8daefdd[23]),
    .b(al_aa3e519e[23]),
    .c(al_ebe24e3d),
    .o({al_c22e023d,al_a972f2b7[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_13acf86f (
    .a(al_f8daefdd[24]),
    .b(al_aa3e519e[24]),
    .c(al_c22e023d),
    .o({al_7aed21eb,al_a972f2b7[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2d4b19b0 (
    .a(al_f8daefdd[25]),
    .b(al_aa3e519e[25]),
    .c(al_7aed21eb),
    .o({al_de434a70,al_a972f2b7[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a26775c (
    .a(al_f8daefdd[26]),
    .b(al_aa3e519e[26]),
    .c(al_de434a70),
    .o({al_4026dc20,al_a972f2b7[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b1c2ed24 (
    .a(al_f8daefdd[27]),
    .b(al_aa3e519e[27]),
    .c(al_4026dc20),
    .o({al_7c090755,al_a972f2b7[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dad5f785 (
    .a(al_f8daefdd[28]),
    .b(al_aa3e519e[28]),
    .c(al_7c090755),
    .o({al_ae7b2873,al_a972f2b7[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b6cb8a97 (
    .a(al_f8daefdd[29]),
    .b(al_aa3e519e[29]),
    .c(al_ae7b2873),
    .o({al_e8aded2c,al_a972f2b7[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b693e974 (
    .a(al_f8daefdd[30]),
    .b(al_aa3e519e[30]),
    .c(al_e8aded2c),
    .o({al_d89660dd,al_a972f2b7[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d2944d0a (
    .a(al_f8daefdd[31]),
    .b(al_aa3e519e[31]),
    .c(al_d89660dd),
    .o({al_a0eacc1c,al_a972f2b7[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dd08739a (
    .a(al_f8daefdd[32]),
    .b(al_aa3e519e[32]),
    .c(al_a0eacc1c),
    .o({al_371958b8,al_a972f2b7[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_744dc21e (
    .a(al_f8daefdd[33]),
    .b(al_aa3e519e[33]),
    .c(al_371958b8),
    .o({al_69ee2d7e,al_a972f2b7[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40b38898 (
    .a(al_f8daefdd[34]),
    .b(al_aa3e519e[34]),
    .c(al_69ee2d7e),
    .o({al_a313220b,al_a972f2b7[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c4e6d5a7 (
    .a(al_f8daefdd[35]),
    .b(al_aa3e519e[35]),
    .c(al_a313220b),
    .o({al_cde03fa5,al_a972f2b7[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ae2a886e (
    .a(al_f8daefdd[36]),
    .b(al_aa3e519e[36]),
    .c(al_cde03fa5),
    .o({al_47e767,al_a972f2b7[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_42e58b6b (
    .a(al_f8daefdd[37]),
    .b(al_aa3e519e[37]),
    .c(al_47e767),
    .o({al_160b1ef,al_a972f2b7[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_da1bd508 (
    .a(al_f8daefdd[38]),
    .b(1'b0),
    .c(al_160b1ef),
    .o({al_8178bce7,open_n178}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6cc5885c (
    .a(1'b0),
    .b(1'b1),
    .c(al_8178bce7),
    .o({open_n179,al_ebc6f995}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_71ab9944 (
    .a(al_f8daefdd[10]),
    .b(al_a972f2b7[4]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_54a67aa9 (
    .a(al_f8daefdd[11]),
    .b(al_a972f2b7[5]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2244d63b (
    .a(al_f8daefdd[12]),
    .b(al_a972f2b7[6]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_18a213a6 (
    .a(al_f8daefdd[13]),
    .b(al_a972f2b7[7]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5666563c (
    .a(al_f8daefdd[14]),
    .b(al_a972f2b7[8]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cbff1c92 (
    .a(al_f8daefdd[15]),
    .b(al_a972f2b7[9]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9d6fcc57 (
    .a(al_f8daefdd[16]),
    .b(al_a972f2b7[10]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a4116e83 (
    .a(al_f8daefdd[17]),
    .b(al_a972f2b7[11]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a50cfc7f (
    .a(al_f8daefdd[18]),
    .b(al_a972f2b7[12]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a3d08383 (
    .a(al_f8daefdd[19]),
    .b(al_a972f2b7[13]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_45a4b403 (
    .a(al_f8daefdd[20]),
    .b(al_a972f2b7[14]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7f1c3f0c (
    .a(al_f8daefdd[21]),
    .b(al_a972f2b7[15]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_aca64528 (
    .a(al_f8daefdd[22]),
    .b(al_a972f2b7[16]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ba3ebd3e (
    .a(al_f8daefdd[23]),
    .b(al_a972f2b7[17]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e1e7a64e (
    .a(al_f8daefdd[24]),
    .b(al_a972f2b7[18]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9c82f114 (
    .a(al_f8daefdd[25]),
    .b(al_a972f2b7[19]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6615d509 (
    .a(al_f8daefdd[26]),
    .b(al_a972f2b7[20]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_243db275 (
    .a(al_f8daefdd[27]),
    .b(al_a972f2b7[21]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c50aea33 (
    .a(al_f8daefdd[28]),
    .b(al_a972f2b7[22]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9bdff1eb (
    .a(al_f8daefdd[29]),
    .b(al_a972f2b7[23]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9c3a20ec (
    .a(al_f8daefdd[30]),
    .b(al_a972f2b7[24]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_572e4896 (
    .a(al_f8daefdd[31]),
    .b(al_a972f2b7[25]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d89319c5 (
    .a(al_f8daefdd[32]),
    .b(al_a972f2b7[26]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_901d36e (
    .a(al_f8daefdd[33]),
    .b(al_a972f2b7[27]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7bc4ae59 (
    .a(al_f8daefdd[34]),
    .b(al_a972f2b7[28]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e0330ff8 (
    .a(al_f8daefdd[35]),
    .b(al_a972f2b7[29]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_35e91380 (
    .a(al_f8daefdd[36]),
    .b(al_a972f2b7[30]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_db56aaf5 (
    .a(al_f8daefdd[37]),
    .b(al_a972f2b7[31]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[37]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3edba449 (
    .a(al_f8daefdd[6]),
    .b(al_a972f2b7[0]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_74cc953 (
    .a(al_f8daefdd[7]),
    .b(al_a972f2b7[1]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a0761a7e (
    .a(al_f8daefdd[8]),
    .b(al_a972f2b7[2]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8cf59845 (
    .a(al_f8daefdd[9]),
    .b(al_a972f2b7[3]),
    .c(al_ebc6f995),
    .o(al_c5d46f6b[9]));
  AL_DFF_X al_293ad1c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8daefdd[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[0]));
  AL_DFF_X al_e273603a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[9]));
  AL_DFF_X al_eb3af9ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[10]));
  AL_DFF_X al_2ab54ae2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[11]));
  AL_DFF_X al_9cdbffbb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[12]));
  AL_DFF_X al_b32f6730 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[13]));
  AL_DFF_X al_101f1373 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[14]));
  AL_DFF_X al_f1cebccb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[15]));
  AL_DFF_X al_ebd82a1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[16]));
  AL_DFF_X al_c4232423 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[17]));
  AL_DFF_X al_97644ffa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[18]));
  AL_DFF_X al_ec6bc5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8daefdd[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[1]));
  AL_DFF_X al_73028f0b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[19]));
  AL_DFF_X al_feeb9917 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[20]));
  AL_DFF_X al_e48ee2a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[21]));
  AL_DFF_X al_f8a4bb5c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[22]));
  AL_DFF_X al_b8abee01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[23]));
  AL_DFF_X al_d6dcbd14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[24]));
  AL_DFF_X al_a8bfbe98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[25]));
  AL_DFF_X al_20a53a7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[26]));
  AL_DFF_X al_4cc27ecc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[27]));
  AL_DFF_X al_1083ddf2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[28]));
  AL_DFF_X al_b9b6c9ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8daefdd[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[2]));
  AL_DFF_X al_40bfdc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[29]));
  AL_DFF_X al_ee747f05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[30]));
  AL_DFF_X al_7c958536 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[31]));
  AL_DFF_X al_20e72348 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[32]));
  AL_DFF_X al_d655c53f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[33]));
  AL_DFF_X al_b8949918 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[34]));
  AL_DFF_X al_7304a692 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[35]));
  AL_DFF_X al_cdd1c3eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[36]));
  AL_DFF_X al_6fa384d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[37]));
  AL_DFF_X al_81225382 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8daefdd[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[3]));
  AL_DFF_X al_71dc030 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8daefdd[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[4]));
  AL_DFF_X al_4f4ee97c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f8daefdd[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[5]));
  AL_DFF_X al_ac7cc553 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[6]));
  AL_DFF_X al_cca77c36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[7]));
  AL_DFF_X al_2286bccb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c5d46f6b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_32798732[8]));
  AL_DFF_X al_5d1598ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ebc6f995),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[0]));
  AL_DFF_X al_32951c92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[9]));
  AL_DFF_X al_39579f65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[10]));
  AL_DFF_X al_16fdf2b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[11]));
  AL_DFF_X al_cf4b63f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[12]));
  AL_DFF_X al_9d3acf92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[13]));
  AL_DFF_X al_a398bfa2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[14]));
  AL_DFF_X al_2e765e3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[15]));
  AL_DFF_X al_625d32bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[16]));
  AL_DFF_X al_c640881b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[17]));
  AL_DFF_X al_5b2e884c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[18]));
  AL_DFF_X al_b5f5773a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[1]));
  AL_DFF_X al_84eae558 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[19]));
  AL_DFF_X al_9e9719f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[20]));
  AL_DFF_X al_917b17fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[21]));
  AL_DFF_X al_802a7988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[22]));
  AL_DFF_X al_ab0b3778 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[23]));
  AL_DFF_X al_7d107297 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[24]));
  AL_DFF_X al_6df64e28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[25]));
  AL_DFF_X al_1d13265f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[26]));
  AL_DFF_X al_aa20d936 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[27]));
  AL_DFF_X al_10ee5f6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[28]));
  AL_DFF_X al_d4b19610 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[2]));
  AL_DFF_X al_5c480a70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[29]));
  AL_DFF_X al_9f413170 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[30]));
  AL_DFF_X al_17a0e5d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[31]));
  AL_DFF_X al_8bcd9c58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[32]));
  AL_DFF_X al_d4f48a16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[33]));
  AL_DFF_X al_faf45239 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[34]));
  AL_DFF_X al_ea147863 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[35]));
  AL_DFF_X al_1e3c7a02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[36]));
  AL_DFF_X al_1f5c3b53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[37]));
  AL_DFF_X al_20b4c236 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[38]));
  AL_DFF_X al_99a6b320 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[3]));
  AL_DFF_X al_1ee487c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[39]));
  AL_DFF_X al_80e6e055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[40]));
  AL_DFF_X al_ecc531ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[41]));
  AL_DFF_X al_b4c42ab2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[4]));
  AL_DFF_X al_2bfb4545 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[5]));
  AL_DFF_X al_e2760c14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[6]));
  AL_DFF_X al_c572e0ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[7]));
  AL_DFF_X al_6b38246c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3357c8f6[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7d914746[8]));
  AL_DFF_X al_6f9934b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_993138f9[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d5d72c9e[0]));
  AL_DFF_X al_fe59b6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[9]));
  AL_DFF_X al_6924e12a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[10]));
  AL_DFF_X al_669f4826 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[11]));
  AL_DFF_X al_41365748 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[12]));
  AL_DFF_X al_185d9f46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[13]));
  AL_DFF_X al_745578bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[14]));
  AL_DFF_X al_7ea6c7a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[15]));
  AL_DFF_X al_48067f15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[16]));
  AL_DFF_X al_fc12f39c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[17]));
  AL_DFF_X al_ced906f2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[18]));
  AL_DFF_X al_9fd700e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[19]));
  AL_DFF_X al_10de2a57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[20]));
  AL_DFF_X al_4b737310 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[21]));
  AL_DFF_X al_5b7ac647 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[22]));
  AL_DFF_X al_5e8f7043 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[23]));
  AL_DFF_X al_419d9dbc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[24]));
  AL_DFF_X al_b60b75e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[25]));
  AL_DFF_X al_98d3f79c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[26]));
  AL_DFF_X al_d5542b6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[27]));
  AL_DFF_X al_66fc636c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[28]));
  AL_DFF_X al_a86bb122 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[29]));
  AL_DFF_X al_9f9daa0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[30]));
  AL_DFF_X al_35deae87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[31]));
  AL_DFF_X al_9b9c8cd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[32]));
  AL_DFF_X al_ef55f399 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[33]));
  AL_DFF_X al_93dff3b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[34]));
  AL_DFF_X al_ae09e20c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[35]));
  AL_DFF_X al_697e7e88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[4]));
  AL_DFF_X al_e16f27ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[5]));
  AL_DFF_X al_c68224a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[6]));
  AL_DFF_X al_afa2bf42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[7]));
  AL_DFF_X al_65ef664f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5e4a13f0[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22838ccb[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_643850ad (
    .a(1'b0),
    .o({al_bc6f54a9,open_n182}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_418ea284 (
    .a(al_32798732[5]),
    .b(al_5e4a13f0[5]),
    .c(al_bc6f54a9),
    .o({al_1a110913,al_a7bae927[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c3dd09e (
    .a(al_32798732[6]),
    .b(al_5e4a13f0[6]),
    .c(al_1a110913),
    .o({al_b4aada3d,al_a7bae927[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9199d8e5 (
    .a(al_32798732[7]),
    .b(al_5e4a13f0[7]),
    .c(al_b4aada3d),
    .o({al_5f7332b4,al_a7bae927[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e85aee19 (
    .a(al_32798732[8]),
    .b(al_5e4a13f0[8]),
    .c(al_5f7332b4),
    .o({al_64d12b15,al_a7bae927[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1aeebf78 (
    .a(al_32798732[9]),
    .b(al_5e4a13f0[9]),
    .c(al_64d12b15),
    .o({al_13e60b1b,al_a7bae927[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c64e068d (
    .a(al_32798732[10]),
    .b(al_5e4a13f0[10]),
    .c(al_13e60b1b),
    .o({al_e0e9a4f3,al_a7bae927[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f35fa265 (
    .a(al_32798732[11]),
    .b(al_5e4a13f0[11]),
    .c(al_e0e9a4f3),
    .o({al_dbf8fa9d,al_a7bae927[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1d624976 (
    .a(al_32798732[12]),
    .b(al_5e4a13f0[12]),
    .c(al_dbf8fa9d),
    .o({al_f5f324f,al_a7bae927[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5f4079c8 (
    .a(al_32798732[13]),
    .b(al_5e4a13f0[13]),
    .c(al_f5f324f),
    .o({al_6766b849,al_a7bae927[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_81d6aa7 (
    .a(al_32798732[14]),
    .b(al_5e4a13f0[14]),
    .c(al_6766b849),
    .o({al_143e4872,al_a7bae927[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b48f4bb (
    .a(al_32798732[15]),
    .b(al_5e4a13f0[15]),
    .c(al_143e4872),
    .o({al_a477b479,al_a7bae927[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a27c8b6a (
    .a(al_32798732[16]),
    .b(al_5e4a13f0[16]),
    .c(al_a477b479),
    .o({al_8bc3354,al_a7bae927[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_90d48ce1 (
    .a(al_32798732[17]),
    .b(al_5e4a13f0[17]),
    .c(al_8bc3354),
    .o({al_1e6bd6a1,al_a7bae927[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d2f1a541 (
    .a(al_32798732[18]),
    .b(al_5e4a13f0[18]),
    .c(al_1e6bd6a1),
    .o({al_e69868df,al_a7bae927[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eb15bee9 (
    .a(al_32798732[19]),
    .b(al_5e4a13f0[19]),
    .c(al_e69868df),
    .o({al_ae74b6ce,al_a7bae927[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9956dcfc (
    .a(al_32798732[20]),
    .b(al_5e4a13f0[20]),
    .c(al_ae74b6ce),
    .o({al_9290634f,al_a7bae927[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3169c5d2 (
    .a(al_32798732[21]),
    .b(al_5e4a13f0[21]),
    .c(al_9290634f),
    .o({al_7af9dc,al_a7bae927[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_74fa5eae (
    .a(al_32798732[22]),
    .b(al_5e4a13f0[22]),
    .c(al_7af9dc),
    .o({al_8084b00c,al_a7bae927[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f732be13 (
    .a(al_32798732[23]),
    .b(al_5e4a13f0[23]),
    .c(al_8084b00c),
    .o({al_b760f405,al_a7bae927[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bbffa5f8 (
    .a(al_32798732[24]),
    .b(al_5e4a13f0[24]),
    .c(al_b760f405),
    .o({al_65d1cfc2,al_a7bae927[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_13b72bf5 (
    .a(al_32798732[25]),
    .b(al_5e4a13f0[25]),
    .c(al_65d1cfc2),
    .o({al_117e7922,al_a7bae927[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a1da72be (
    .a(al_32798732[26]),
    .b(al_5e4a13f0[26]),
    .c(al_117e7922),
    .o({al_633d0b30,al_a7bae927[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a5cf647 (
    .a(al_32798732[27]),
    .b(al_5e4a13f0[27]),
    .c(al_633d0b30),
    .o({al_b3570833,al_a7bae927[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2fb8dfd8 (
    .a(al_32798732[28]),
    .b(al_5e4a13f0[28]),
    .c(al_b3570833),
    .o({al_b9b8f3e1,al_a7bae927[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d8df4ae7 (
    .a(al_32798732[29]),
    .b(al_5e4a13f0[29]),
    .c(al_b9b8f3e1),
    .o({al_37f2f859,al_a7bae927[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_54bb3efd (
    .a(al_32798732[30]),
    .b(al_5e4a13f0[30]),
    .c(al_37f2f859),
    .o({al_691ab75e,al_a7bae927[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9e84b6a9 (
    .a(al_32798732[31]),
    .b(al_5e4a13f0[31]),
    .c(al_691ab75e),
    .o({al_78df4457,al_a7bae927[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e964dfed (
    .a(al_32798732[32]),
    .b(al_5e4a13f0[32]),
    .c(al_78df4457),
    .o({al_ea3d8437,al_a7bae927[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2f68adfc (
    .a(al_32798732[33]),
    .b(al_5e4a13f0[33]),
    .c(al_ea3d8437),
    .o({al_d03ec855,al_a7bae927[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a67bd437 (
    .a(al_32798732[34]),
    .b(al_5e4a13f0[34]),
    .c(al_d03ec855),
    .o({al_d1805774,al_a7bae927[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4f625637 (
    .a(al_32798732[35]),
    .b(al_5e4a13f0[35]),
    .c(al_d1805774),
    .o({al_b2501f7c,al_a7bae927[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6775e7e0 (
    .a(al_32798732[36]),
    .b(al_5e4a13f0[36]),
    .c(al_b2501f7c),
    .o({al_2e361070,al_a7bae927[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_15253c25 (
    .a(al_32798732[37]),
    .b(1'b0),
    .c(al_2e361070),
    .o({al_9b14b36d,open_n183}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_835bdb60 (
    .a(1'b0),
    .b(1'b1),
    .c(al_9b14b36d),
    .o({open_n184,al_e0fb24bc}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_da078be (
    .a(al_32798732[10]),
    .b(al_a7bae927[5]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2265d26a (
    .a(al_32798732[11]),
    .b(al_a7bae927[6]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fa5777f3 (
    .a(al_32798732[12]),
    .b(al_a7bae927[7]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_19e07f88 (
    .a(al_32798732[13]),
    .b(al_a7bae927[8]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3b75f218 (
    .a(al_32798732[14]),
    .b(al_a7bae927[9]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3265ba00 (
    .a(al_32798732[15]),
    .b(al_a7bae927[10]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6e17e85a (
    .a(al_32798732[16]),
    .b(al_a7bae927[11]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f22ed44 (
    .a(al_32798732[17]),
    .b(al_a7bae927[12]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2032c4cd (
    .a(al_32798732[18]),
    .b(al_a7bae927[13]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_dda949eb (
    .a(al_32798732[19]),
    .b(al_a7bae927[14]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_293248fb (
    .a(al_32798732[20]),
    .b(al_a7bae927[15]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_580ba467 (
    .a(al_32798732[21]),
    .b(al_a7bae927[16]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ecc4bb7 (
    .a(al_32798732[22]),
    .b(al_a7bae927[17]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8a4dc70d (
    .a(al_32798732[23]),
    .b(al_a7bae927[18]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d7a0c6a9 (
    .a(al_32798732[24]),
    .b(al_a7bae927[19]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4c92c3ee (
    .a(al_32798732[25]),
    .b(al_a7bae927[20]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f35f5021 (
    .a(al_32798732[26]),
    .b(al_a7bae927[21]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a4be692a (
    .a(al_32798732[27]),
    .b(al_a7bae927[22]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f94c1fb8 (
    .a(al_32798732[28]),
    .b(al_a7bae927[23]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8bedc32e (
    .a(al_32798732[29]),
    .b(al_a7bae927[24]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_28f3a232 (
    .a(al_32798732[30]),
    .b(al_a7bae927[25]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_67208cda (
    .a(al_32798732[31]),
    .b(al_a7bae927[26]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5886a5e2 (
    .a(al_32798732[32]),
    .b(al_a7bae927[27]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bd0e50e6 (
    .a(al_32798732[33]),
    .b(al_a7bae927[28]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b24ef160 (
    .a(al_32798732[34]),
    .b(al_a7bae927[29]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bfac3161 (
    .a(al_32798732[35]),
    .b(al_a7bae927[30]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f501dab3 (
    .a(al_32798732[36]),
    .b(al_a7bae927[31]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[36]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_116eb862 (
    .a(al_32798732[5]),
    .b(al_a7bae927[0]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_755c9ba8 (
    .a(al_32798732[6]),
    .b(al_a7bae927[1]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d59a5af6 (
    .a(al_32798732[7]),
    .b(al_a7bae927[2]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_dfdce7fd (
    .a(al_32798732[8]),
    .b(al_a7bae927[3]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a07bbfa6 (
    .a(al_32798732[9]),
    .b(al_a7bae927[4]),
    .c(al_e0fb24bc),
    .o(al_93803eaa[9]));
  AL_DFF_X al_4708dc04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32798732[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[0]));
  AL_DFF_X al_ac85863 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[9]));
  AL_DFF_X al_ca2c8b85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[10]));
  AL_DFF_X al_5bca3799 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[11]));
  AL_DFF_X al_904698a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[12]));
  AL_DFF_X al_5ebc0a69 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[13]));
  AL_DFF_X al_5f495942 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[14]));
  AL_DFF_X al_d028f683 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[15]));
  AL_DFF_X al_7c70e235 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[16]));
  AL_DFF_X al_b4e776d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[17]));
  AL_DFF_X al_b9727a83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[18]));
  AL_DFF_X al_97938a63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32798732[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[1]));
  AL_DFF_X al_7a5f8d79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[19]));
  AL_DFF_X al_fd451f8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[20]));
  AL_DFF_X al_d0d8eebd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[21]));
  AL_DFF_X al_a2c9bac7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[22]));
  AL_DFF_X al_73ce48c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[23]));
  AL_DFF_X al_b5ce15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[24]));
  AL_DFF_X al_b2d1969c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[25]));
  AL_DFF_X al_ce5fc42d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[26]));
  AL_DFF_X al_fc9bd65c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[27]));
  AL_DFF_X al_b033aacc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[28]));
  AL_DFF_X al_e2e70869 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32798732[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[2]));
  AL_DFF_X al_bcb9058 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[29]));
  AL_DFF_X al_bcea9ffc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[30]));
  AL_DFF_X al_cd9594ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[31]));
  AL_DFF_X al_779acff7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[32]));
  AL_DFF_X al_b946209c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[33]));
  AL_DFF_X al_be5fb5fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[34]));
  AL_DFF_X al_9bcb5111 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[35]));
  AL_DFF_X al_3607f476 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[36]));
  AL_DFF_X al_ab306ec1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32798732[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[3]));
  AL_DFF_X al_78eca474 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_32798732[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[4]));
  AL_DFF_X al_c7ca66a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[5]));
  AL_DFF_X al_b9639eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[6]));
  AL_DFF_X al_dfebb648 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[7]));
  AL_DFF_X al_5efd22aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_93803eaa[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2f60c4e5[8]));
  AL_DFF_X al_da1f400d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_e0fb24bc),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[0]));
  AL_DFF_X al_65d26122 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[9]));
  AL_DFF_X al_8a789ec0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[10]));
  AL_DFF_X al_6d999a2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[11]));
  AL_DFF_X al_20788507 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[12]));
  AL_DFF_X al_f31b7af1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[13]));
  AL_DFF_X al_b60cf355 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[14]));
  AL_DFF_X al_74c7d9a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[15]));
  AL_DFF_X al_991c4e2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[16]));
  AL_DFF_X al_5588f879 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[17]));
  AL_DFF_X al_8ea663a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[18]));
  AL_DFF_X al_74338644 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[1]));
  AL_DFF_X al_e09e0f98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[19]));
  AL_DFF_X al_9b7dd49f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[20]));
  AL_DFF_X al_9a92b267 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[21]));
  AL_DFF_X al_8a58cf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[22]));
  AL_DFF_X al_dbfb5e54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[23]));
  AL_DFF_X al_259b7673 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[24]));
  AL_DFF_X al_fd91326c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[25]));
  AL_DFF_X al_9991d428 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[26]));
  AL_DFF_X al_65728ce2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[27]));
  AL_DFF_X al_6ecb581f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[28]));
  AL_DFF_X al_374bc0b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[2]));
  AL_DFF_X al_462032d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[29]));
  AL_DFF_X al_54a56d9e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[30]));
  AL_DFF_X al_a169dba1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[31]));
  AL_DFF_X al_72fa9f96 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[32]));
  AL_DFF_X al_49eadba7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[33]));
  AL_DFF_X al_da9a624 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[34]));
  AL_DFF_X al_c25a5b6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[35]));
  AL_DFF_X al_d4907dfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[36]));
  AL_DFF_X al_bfa4f64c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[37]));
  AL_DFF_X al_7202fc5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[38]));
  AL_DFF_X al_b78fb002 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[3]));
  AL_DFF_X al_a7e2fa27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[39]));
  AL_DFF_X al_e215ea76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[40]));
  AL_DFF_X al_749c4d3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[41]));
  AL_DFF_X al_2d9562ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[42]));
  AL_DFF_X al_1cd1d84b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[4]));
  AL_DFF_X al_197a56f7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[5]));
  AL_DFF_X al_d42a821d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[6]));
  AL_DFF_X al_3d0c7160 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[7]));
  AL_DFF_X al_dcddaad5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d914746[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_97fb94a7[8]));
  AL_DFF_X al_cdb462fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d5d72c9e[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2be1e26f[0]));
  AL_DFF_X al_d5b032d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[9]));
  AL_DFF_X al_deadec6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[10]));
  AL_DFF_X al_9eea0eac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[11]));
  AL_DFF_X al_59716c0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[12]));
  AL_DFF_X al_952cb9eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[13]));
  AL_DFF_X al_57f0b32e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[14]));
  AL_DFF_X al_bf84f76c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[15]));
  AL_DFF_X al_2a359e4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[16]));
  AL_DFF_X al_760fa473 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[17]));
  AL_DFF_X al_84310019 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[18]));
  AL_DFF_X al_c2af3d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[19]));
  AL_DFF_X al_f9f76313 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[20]));
  AL_DFF_X al_4f1a9ad3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[21]));
  AL_DFF_X al_384e9fa6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[22]));
  AL_DFF_X al_fab68763 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[23]));
  AL_DFF_X al_44fa19bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[24]));
  AL_DFF_X al_a26f7810 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[25]));
  AL_DFF_X al_914562d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[26]));
  AL_DFF_X al_e518bc9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[27]));
  AL_DFF_X al_59b83495 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[28]));
  AL_DFF_X al_7ed9a817 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[29]));
  AL_DFF_X al_bd3fdca4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[30]));
  AL_DFF_X al_47770b5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[31]));
  AL_DFF_X al_c3bbd594 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[32]));
  AL_DFF_X al_3f42476c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[33]));
  AL_DFF_X al_c512e94c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[34]));
  AL_DFF_X al_be101c6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[3]));
  AL_DFF_X al_957b9174 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[4]));
  AL_DFF_X al_1da77d24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[5]));
  AL_DFF_X al_2c193140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[6]));
  AL_DFF_X al_a2c23377 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[7]));
  AL_DFF_X al_62741d15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22838ccb[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_44122f34[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_47a60b4b (
    .a(1'b0),
    .o({al_2434069f,open_n187}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_92b009a0 (
    .a(al_2f60c4e5[4]),
    .b(al_22838ccb[4]),
    .c(al_2434069f),
    .o({al_f06b68e,al_6c10dd8f[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8f11539d (
    .a(al_2f60c4e5[5]),
    .b(al_22838ccb[5]),
    .c(al_f06b68e),
    .o({al_eed0f9b1,al_6c10dd8f[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_43e0913e (
    .a(al_2f60c4e5[6]),
    .b(al_22838ccb[6]),
    .c(al_eed0f9b1),
    .o({al_3fdcd506,al_6c10dd8f[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f599d8b5 (
    .a(al_2f60c4e5[7]),
    .b(al_22838ccb[7]),
    .c(al_3fdcd506),
    .o({al_8b101552,al_6c10dd8f[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7d1bdff9 (
    .a(al_2f60c4e5[8]),
    .b(al_22838ccb[8]),
    .c(al_8b101552),
    .o({al_6d93b728,al_6c10dd8f[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cba1d9a8 (
    .a(al_2f60c4e5[9]),
    .b(al_22838ccb[9]),
    .c(al_6d93b728),
    .o({al_fef237c0,al_6c10dd8f[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e2d095a1 (
    .a(al_2f60c4e5[10]),
    .b(al_22838ccb[10]),
    .c(al_fef237c0),
    .o({al_1a734e00,al_6c10dd8f[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_99733a6c (
    .a(al_2f60c4e5[11]),
    .b(al_22838ccb[11]),
    .c(al_1a734e00),
    .o({al_450062f6,al_6c10dd8f[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bf982d41 (
    .a(al_2f60c4e5[12]),
    .b(al_22838ccb[12]),
    .c(al_450062f6),
    .o({al_96c7325f,al_6c10dd8f[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f6f3f823 (
    .a(al_2f60c4e5[13]),
    .b(al_22838ccb[13]),
    .c(al_96c7325f),
    .o({al_34dcc703,al_6c10dd8f[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a9e8f4d3 (
    .a(al_2f60c4e5[14]),
    .b(al_22838ccb[14]),
    .c(al_34dcc703),
    .o({al_8581252c,al_6c10dd8f[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_39ce2927 (
    .a(al_2f60c4e5[15]),
    .b(al_22838ccb[15]),
    .c(al_8581252c),
    .o({al_47ef5621,al_6c10dd8f[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3abfb75f (
    .a(al_2f60c4e5[16]),
    .b(al_22838ccb[16]),
    .c(al_47ef5621),
    .o({al_5595f015,al_6c10dd8f[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e7207588 (
    .a(al_2f60c4e5[17]),
    .b(al_22838ccb[17]),
    .c(al_5595f015),
    .o({al_7cd1dfe0,al_6c10dd8f[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_998f10f7 (
    .a(al_2f60c4e5[18]),
    .b(al_22838ccb[18]),
    .c(al_7cd1dfe0),
    .o({al_3baab685,al_6c10dd8f[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1892320d (
    .a(al_2f60c4e5[19]),
    .b(al_22838ccb[19]),
    .c(al_3baab685),
    .o({al_bfe04e37,al_6c10dd8f[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_280a623f (
    .a(al_2f60c4e5[20]),
    .b(al_22838ccb[20]),
    .c(al_bfe04e37),
    .o({al_ff7baa95,al_6c10dd8f[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2b39956 (
    .a(al_2f60c4e5[21]),
    .b(al_22838ccb[21]),
    .c(al_ff7baa95),
    .o({al_4beff26f,al_6c10dd8f[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b0a85acd (
    .a(al_2f60c4e5[22]),
    .b(al_22838ccb[22]),
    .c(al_4beff26f),
    .o({al_215503f7,al_6c10dd8f[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5ed0308e (
    .a(al_2f60c4e5[23]),
    .b(al_22838ccb[23]),
    .c(al_215503f7),
    .o({al_6ebcb190,al_6c10dd8f[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a63c1d0b (
    .a(al_2f60c4e5[24]),
    .b(al_22838ccb[24]),
    .c(al_6ebcb190),
    .o({al_e3b23b3d,al_6c10dd8f[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_abb69b5d (
    .a(al_2f60c4e5[25]),
    .b(al_22838ccb[25]),
    .c(al_e3b23b3d),
    .o({al_27782d3b,al_6c10dd8f[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b3ce804b (
    .a(al_2f60c4e5[26]),
    .b(al_22838ccb[26]),
    .c(al_27782d3b),
    .o({al_96a09b29,al_6c10dd8f[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_52edbe09 (
    .a(al_2f60c4e5[27]),
    .b(al_22838ccb[27]),
    .c(al_96a09b29),
    .o({al_f5c79977,al_6c10dd8f[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a86aa0e7 (
    .a(al_2f60c4e5[28]),
    .b(al_22838ccb[28]),
    .c(al_f5c79977),
    .o({al_d0973a8a,al_6c10dd8f[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9da9b731 (
    .a(al_2f60c4e5[29]),
    .b(al_22838ccb[29]),
    .c(al_d0973a8a),
    .o({al_53ed7af5,al_6c10dd8f[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_56f58d92 (
    .a(al_2f60c4e5[30]),
    .b(al_22838ccb[30]),
    .c(al_53ed7af5),
    .o({al_f5a1ca8f,al_6c10dd8f[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_24d8384d (
    .a(al_2f60c4e5[31]),
    .b(al_22838ccb[31]),
    .c(al_f5a1ca8f),
    .o({al_c40e7d13,al_6c10dd8f[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_53d089f7 (
    .a(al_2f60c4e5[32]),
    .b(al_22838ccb[32]),
    .c(al_c40e7d13),
    .o({al_b434c7b1,al_6c10dd8f[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7422e5dc (
    .a(al_2f60c4e5[33]),
    .b(al_22838ccb[33]),
    .c(al_b434c7b1),
    .o({al_8d68d680,al_6c10dd8f[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_869eb0f7 (
    .a(al_2f60c4e5[34]),
    .b(al_22838ccb[34]),
    .c(al_8d68d680),
    .o({al_af211502,al_6c10dd8f[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_cc2795ac (
    .a(al_2f60c4e5[35]),
    .b(al_22838ccb[35]),
    .c(al_af211502),
    .o({al_7b9dbd92,al_6c10dd8f[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bf24850e (
    .a(al_2f60c4e5[36]),
    .b(1'b0),
    .c(al_7b9dbd92),
    .o({al_ce16dbbf,open_n188}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5b9bffc9 (
    .a(1'b0),
    .b(1'b1),
    .c(al_ce16dbbf),
    .o({open_n189,al_95f16875}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f73bac05 (
    .a(al_2f60c4e5[10]),
    .b(al_6c10dd8f[6]),
    .c(al_95f16875),
    .o(al_1a0e1c89[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3512e9c9 (
    .a(al_2f60c4e5[11]),
    .b(al_6c10dd8f[7]),
    .c(al_95f16875),
    .o(al_1a0e1c89[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a1511ea1 (
    .a(al_2f60c4e5[12]),
    .b(al_6c10dd8f[8]),
    .c(al_95f16875),
    .o(al_1a0e1c89[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_341d49c6 (
    .a(al_2f60c4e5[13]),
    .b(al_6c10dd8f[9]),
    .c(al_95f16875),
    .o(al_1a0e1c89[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_34c17589 (
    .a(al_2f60c4e5[14]),
    .b(al_6c10dd8f[10]),
    .c(al_95f16875),
    .o(al_1a0e1c89[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1b845000 (
    .a(al_2f60c4e5[15]),
    .b(al_6c10dd8f[11]),
    .c(al_95f16875),
    .o(al_1a0e1c89[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_be17fb56 (
    .a(al_2f60c4e5[16]),
    .b(al_6c10dd8f[12]),
    .c(al_95f16875),
    .o(al_1a0e1c89[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_414f5dcf (
    .a(al_2f60c4e5[17]),
    .b(al_6c10dd8f[13]),
    .c(al_95f16875),
    .o(al_1a0e1c89[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_28583a07 (
    .a(al_2f60c4e5[18]),
    .b(al_6c10dd8f[14]),
    .c(al_95f16875),
    .o(al_1a0e1c89[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_dfba5d68 (
    .a(al_2f60c4e5[19]),
    .b(al_6c10dd8f[15]),
    .c(al_95f16875),
    .o(al_1a0e1c89[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_db1d6d7e (
    .a(al_2f60c4e5[20]),
    .b(al_6c10dd8f[16]),
    .c(al_95f16875),
    .o(al_1a0e1c89[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c0ec24d2 (
    .a(al_2f60c4e5[21]),
    .b(al_6c10dd8f[17]),
    .c(al_95f16875),
    .o(al_1a0e1c89[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_abf1c561 (
    .a(al_2f60c4e5[22]),
    .b(al_6c10dd8f[18]),
    .c(al_95f16875),
    .o(al_1a0e1c89[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1a1c83f2 (
    .a(al_2f60c4e5[23]),
    .b(al_6c10dd8f[19]),
    .c(al_95f16875),
    .o(al_1a0e1c89[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7095f212 (
    .a(al_2f60c4e5[24]),
    .b(al_6c10dd8f[20]),
    .c(al_95f16875),
    .o(al_1a0e1c89[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8f4d0bd7 (
    .a(al_2f60c4e5[25]),
    .b(al_6c10dd8f[21]),
    .c(al_95f16875),
    .o(al_1a0e1c89[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_37ffa4e3 (
    .a(al_2f60c4e5[26]),
    .b(al_6c10dd8f[22]),
    .c(al_95f16875),
    .o(al_1a0e1c89[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e457d4a8 (
    .a(al_2f60c4e5[27]),
    .b(al_6c10dd8f[23]),
    .c(al_95f16875),
    .o(al_1a0e1c89[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c6b12772 (
    .a(al_2f60c4e5[28]),
    .b(al_6c10dd8f[24]),
    .c(al_95f16875),
    .o(al_1a0e1c89[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bd68d617 (
    .a(al_2f60c4e5[29]),
    .b(al_6c10dd8f[25]),
    .c(al_95f16875),
    .o(al_1a0e1c89[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_577e98ae (
    .a(al_2f60c4e5[30]),
    .b(al_6c10dd8f[26]),
    .c(al_95f16875),
    .o(al_1a0e1c89[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_11bc4312 (
    .a(al_2f60c4e5[31]),
    .b(al_6c10dd8f[27]),
    .c(al_95f16875),
    .o(al_1a0e1c89[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2620103e (
    .a(al_2f60c4e5[32]),
    .b(al_6c10dd8f[28]),
    .c(al_95f16875),
    .o(al_1a0e1c89[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d295ffb0 (
    .a(al_2f60c4e5[33]),
    .b(al_6c10dd8f[29]),
    .c(al_95f16875),
    .o(al_1a0e1c89[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b9488f17 (
    .a(al_2f60c4e5[34]),
    .b(al_6c10dd8f[30]),
    .c(al_95f16875),
    .o(al_1a0e1c89[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d6b70ae3 (
    .a(al_2f60c4e5[35]),
    .b(al_6c10dd8f[31]),
    .c(al_95f16875),
    .o(al_1a0e1c89[35]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ba046516 (
    .a(al_2f60c4e5[4]),
    .b(al_6c10dd8f[0]),
    .c(al_95f16875),
    .o(al_1a0e1c89[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7f669699 (
    .a(al_2f60c4e5[5]),
    .b(al_6c10dd8f[1]),
    .c(al_95f16875),
    .o(al_1a0e1c89[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_62601890 (
    .a(al_2f60c4e5[6]),
    .b(al_6c10dd8f[2]),
    .c(al_95f16875),
    .o(al_1a0e1c89[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8fc93ea (
    .a(al_2f60c4e5[7]),
    .b(al_6c10dd8f[3]),
    .c(al_95f16875),
    .o(al_1a0e1c89[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5630b1cd (
    .a(al_2f60c4e5[8]),
    .b(al_6c10dd8f[4]),
    .c(al_95f16875),
    .o(al_1a0e1c89[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f1ed0315 (
    .a(al_2f60c4e5[9]),
    .b(al_6c10dd8f[5]),
    .c(al_95f16875),
    .o(al_1a0e1c89[9]));
  AL_DFF_X al_297e33ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2f60c4e5[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[0]));
  AL_DFF_X al_4d4a08a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[9]));
  AL_DFF_X al_b1ab8226 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[10]));
  AL_DFF_X al_c8706a59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[11]));
  AL_DFF_X al_3ee62650 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[12]));
  AL_DFF_X al_f2a7217d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[13]));
  AL_DFF_X al_2ccb6358 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[14]));
  AL_DFF_X al_c3064e58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[15]));
  AL_DFF_X al_4e6343cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[16]));
  AL_DFF_X al_429ef820 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[17]));
  AL_DFF_X al_a424b5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[18]));
  AL_DFF_X al_6cfafef6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2f60c4e5[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[1]));
  AL_DFF_X al_32533e28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[19]));
  AL_DFF_X al_925fd8b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[20]));
  AL_DFF_X al_b33e250f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[21]));
  AL_DFF_X al_da7a87be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[22]));
  AL_DFF_X al_ce17b57f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[23]));
  AL_DFF_X al_fe6d33cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[24]));
  AL_DFF_X al_e8d1f36b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[25]));
  AL_DFF_X al_d6ade4a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[26]));
  AL_DFF_X al_6fea30d5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[27]));
  AL_DFF_X al_b04e5be0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[28]));
  AL_DFF_X al_b3ab6e94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2f60c4e5[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[2]));
  AL_DFF_X al_325d4f85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[29]));
  AL_DFF_X al_b48449f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[30]));
  AL_DFF_X al_80c78da5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[31]));
  AL_DFF_X al_4c5e891a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[32]));
  AL_DFF_X al_acdfe54f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[33]));
  AL_DFF_X al_63406e85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[34]));
  AL_DFF_X al_99f1dd6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[35]));
  AL_DFF_X al_85161811 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2f60c4e5[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[3]));
  AL_DFF_X al_9340fccb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[4]));
  AL_DFF_X al_82dfb21e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[5]));
  AL_DFF_X al_152480f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[6]));
  AL_DFF_X al_9d2f4204 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[7]));
  AL_DFF_X al_c9823d8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1a0e1c89[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_167f3ebe[8]));
  AL_DFF_X al_9889ee62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_95f16875),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[0]));
  AL_DFF_X al_8f2b88c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[9]));
  AL_DFF_X al_2e557e98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[10]));
  AL_DFF_X al_7d0a75e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[11]));
  AL_DFF_X al_dc76cb24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[12]));
  AL_DFF_X al_87bb7f95 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[13]));
  AL_DFF_X al_c7af0b5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[14]));
  AL_DFF_X al_53a9eab7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[15]));
  AL_DFF_X al_642cfed9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[16]));
  AL_DFF_X al_84cb943 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[17]));
  AL_DFF_X al_960b5877 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[18]));
  AL_DFF_X al_256c91c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[1]));
  AL_DFF_X al_591a7d1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[19]));
  AL_DFF_X al_8621150e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[20]));
  AL_DFF_X al_7b6c77e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[21]));
  AL_DFF_X al_e572cedd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[22]));
  AL_DFF_X al_46c597ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[23]));
  AL_DFF_X al_b1f5a1e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[24]));
  AL_DFF_X al_77591ddf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[25]));
  AL_DFF_X al_2a33086b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[26]));
  AL_DFF_X al_847fdf73 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[27]));
  AL_DFF_X al_3d0a1d00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[28]));
  AL_DFF_X al_5727194c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[2]));
  AL_DFF_X al_d03f7b0d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[29]));
  AL_DFF_X al_fd9cff98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[30]));
  AL_DFF_X al_f3c9503d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[31]));
  AL_DFF_X al_39e4787d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[32]));
  AL_DFF_X al_b4875ef2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[33]));
  AL_DFF_X al_5f3b4348 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[34]));
  AL_DFF_X al_4f256670 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[35]));
  AL_DFF_X al_ed3bbe93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[36]));
  AL_DFF_X al_f4f8f318 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[37]));
  AL_DFF_X al_819bcb99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[38]));
  AL_DFF_X al_3b54b62d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[3]));
  AL_DFF_X al_f3f742c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[39]));
  AL_DFF_X al_ecf74756 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[40]));
  AL_DFF_X al_8e05e96e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[41]));
  AL_DFF_X al_a2a6562d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[42]));
  AL_DFF_X al_33713275 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[43]));
  AL_DFF_X al_462d5d90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[4]));
  AL_DFF_X al_a668fdf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[5]));
  AL_DFF_X al_400b797f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[6]));
  AL_DFF_X al_706b016c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[7]));
  AL_DFF_X al_5755f6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_97fb94a7[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c2cdf2f1[8]));
  AL_DFF_X al_1b861c7c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2be1e26f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5d2b923b[0]));
  AL_DFF_X al_9db8ebfa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[9]));
  AL_DFF_X al_8c8284d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[10]));
  AL_DFF_X al_4d1f69b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[11]));
  AL_DFF_X al_acc32d4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[12]));
  AL_DFF_X al_d5fc469f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[13]));
  AL_DFF_X al_69d657b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[14]));
  AL_DFF_X al_80b08e18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[15]));
  AL_DFF_X al_836549ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[16]));
  AL_DFF_X al_1241d6c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[17]));
  AL_DFF_X al_779c754 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[18]));
  AL_DFF_X al_348b5d6d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[19]));
  AL_DFF_X al_1f61ae51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[20]));
  AL_DFF_X al_aa028254 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[21]));
  AL_DFF_X al_30af4ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[22]));
  AL_DFF_X al_e754ce3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[23]));
  AL_DFF_X al_84e9b99e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[24]));
  AL_DFF_X al_bef8242c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[25]));
  AL_DFF_X al_54bd11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[26]));
  AL_DFF_X al_4661079e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[27]));
  AL_DFF_X al_e1f82c42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[28]));
  AL_DFF_X al_1ef6d161 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[2]));
  AL_DFF_X al_b3f48cf2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[29]));
  AL_DFF_X al_eb1b2110 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[30]));
  AL_DFF_X al_6a841e4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[31]));
  AL_DFF_X al_13a86e0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[32]));
  AL_DFF_X al_b8624518 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[33]));
  AL_DFF_X al_c911812b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[3]));
  AL_DFF_X al_74b4dfac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[4]));
  AL_DFF_X al_1a978d08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[5]));
  AL_DFF_X al_af2ee180 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[6]));
  AL_DFF_X al_59603df5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[7]));
  AL_DFF_X al_41b1530a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_44122f34[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7e0865ed[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_25d423bb (
    .a(1'b0),
    .o({al_81bff2a0,open_n192}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d923970b (
    .a(al_167f3ebe[3]),
    .b(al_44122f34[3]),
    .c(al_81bff2a0),
    .o({al_b661fbd8,al_a352434c[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e2e605af (
    .a(al_167f3ebe[4]),
    .b(al_44122f34[4]),
    .c(al_b661fbd8),
    .o({al_d0b214a9,al_a352434c[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4dfa71ee (
    .a(al_167f3ebe[5]),
    .b(al_44122f34[5]),
    .c(al_d0b214a9),
    .o({al_9fb02266,al_a352434c[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2454b091 (
    .a(al_167f3ebe[6]),
    .b(al_44122f34[6]),
    .c(al_9fb02266),
    .o({al_c2f2105d,al_a352434c[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c9e2d284 (
    .a(al_167f3ebe[7]),
    .b(al_44122f34[7]),
    .c(al_c2f2105d),
    .o({al_df257acd,al_a352434c[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bd6f50e9 (
    .a(al_167f3ebe[8]),
    .b(al_44122f34[8]),
    .c(al_df257acd),
    .o({al_ceac5249,al_a352434c[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_163d62cc (
    .a(al_167f3ebe[9]),
    .b(al_44122f34[9]),
    .c(al_ceac5249),
    .o({al_a09d4af8,al_a352434c[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7a9d05ae (
    .a(al_167f3ebe[10]),
    .b(al_44122f34[10]),
    .c(al_a09d4af8),
    .o({al_8b2f2894,al_a352434c[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_65d7e508 (
    .a(al_167f3ebe[11]),
    .b(al_44122f34[11]),
    .c(al_8b2f2894),
    .o({al_7ae76686,al_a352434c[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2ea343ec (
    .a(al_167f3ebe[12]),
    .b(al_44122f34[12]),
    .c(al_7ae76686),
    .o({al_4d2bf11f,al_a352434c[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_51a47154 (
    .a(al_167f3ebe[13]),
    .b(al_44122f34[13]),
    .c(al_4d2bf11f),
    .o({al_cedf3c10,al_a352434c[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_190ca347 (
    .a(al_167f3ebe[14]),
    .b(al_44122f34[14]),
    .c(al_cedf3c10),
    .o({al_4e77bfa,al_a352434c[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_25f8000d (
    .a(al_167f3ebe[15]),
    .b(al_44122f34[15]),
    .c(al_4e77bfa),
    .o({al_5efe66e3,al_a352434c[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_222a33ba (
    .a(al_167f3ebe[16]),
    .b(al_44122f34[16]),
    .c(al_5efe66e3),
    .o({al_693c6c75,al_a352434c[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e375bc26 (
    .a(al_167f3ebe[17]),
    .b(al_44122f34[17]),
    .c(al_693c6c75),
    .o({al_822e59ab,al_a352434c[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e8ca130b (
    .a(al_167f3ebe[18]),
    .b(al_44122f34[18]),
    .c(al_822e59ab),
    .o({al_5db6e161,al_a352434c[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_67974ea1 (
    .a(al_167f3ebe[19]),
    .b(al_44122f34[19]),
    .c(al_5db6e161),
    .o({al_34b35b3f,al_a352434c[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_581f19ab (
    .a(al_167f3ebe[20]),
    .b(al_44122f34[20]),
    .c(al_34b35b3f),
    .o({al_5010b887,al_a352434c[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_998f50ce (
    .a(al_167f3ebe[21]),
    .b(al_44122f34[21]),
    .c(al_5010b887),
    .o({al_7d8a00ee,al_a352434c[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_528cfcfa (
    .a(al_167f3ebe[22]),
    .b(al_44122f34[22]),
    .c(al_7d8a00ee),
    .o({al_9bd13530,al_a352434c[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b5809f57 (
    .a(al_167f3ebe[23]),
    .b(al_44122f34[23]),
    .c(al_9bd13530),
    .o({al_a0c66e60,al_a352434c[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_729666d (
    .a(al_167f3ebe[24]),
    .b(al_44122f34[24]),
    .c(al_a0c66e60),
    .o({al_aab46c70,al_a352434c[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_54c3db77 (
    .a(al_167f3ebe[25]),
    .b(al_44122f34[25]),
    .c(al_aab46c70),
    .o({al_7b742de5,al_a352434c[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_23172368 (
    .a(al_167f3ebe[26]),
    .b(al_44122f34[26]),
    .c(al_7b742de5),
    .o({al_5b895c4d,al_a352434c[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_aaa06ecf (
    .a(al_167f3ebe[27]),
    .b(al_44122f34[27]),
    .c(al_5b895c4d),
    .o({al_8526f7d0,al_a352434c[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_43b186df (
    .a(al_167f3ebe[28]),
    .b(al_44122f34[28]),
    .c(al_8526f7d0),
    .o({al_3dd7b884,al_a352434c[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_eda07b06 (
    .a(al_167f3ebe[29]),
    .b(al_44122f34[29]),
    .c(al_3dd7b884),
    .o({al_9c8e7269,al_a352434c[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_976ab2f7 (
    .a(al_167f3ebe[30]),
    .b(al_44122f34[30]),
    .c(al_9c8e7269),
    .o({al_216fbee,al_a352434c[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3164c173 (
    .a(al_167f3ebe[31]),
    .b(al_44122f34[31]),
    .c(al_216fbee),
    .o({al_fdd42739,al_a352434c[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5c892736 (
    .a(al_167f3ebe[32]),
    .b(al_44122f34[32]),
    .c(al_fdd42739),
    .o({al_ed1e8e02,al_a352434c[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_338db74e (
    .a(al_167f3ebe[33]),
    .b(al_44122f34[33]),
    .c(al_ed1e8e02),
    .o({al_8208c979,al_a352434c[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_23bdac46 (
    .a(al_167f3ebe[34]),
    .b(al_44122f34[34]),
    .c(al_8208c979),
    .o({al_2842b1a1,al_a352434c[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4b6453b1 (
    .a(al_167f3ebe[35]),
    .b(1'b0),
    .c(al_2842b1a1),
    .o({al_594d587,open_n193}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_18fae787 (
    .a(1'b0),
    .b(1'b1),
    .c(al_594d587),
    .o({open_n194,al_f57392c}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4ba128b3 (
    .a(al_167f3ebe[10]),
    .b(al_a352434c[7]),
    .c(al_f57392c),
    .o(al_7452903f[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4766c47a (
    .a(al_167f3ebe[11]),
    .b(al_a352434c[8]),
    .c(al_f57392c),
    .o(al_7452903f[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_516ad1a6 (
    .a(al_167f3ebe[12]),
    .b(al_a352434c[9]),
    .c(al_f57392c),
    .o(al_7452903f[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_82c7ca23 (
    .a(al_167f3ebe[13]),
    .b(al_a352434c[10]),
    .c(al_f57392c),
    .o(al_7452903f[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f094c918 (
    .a(al_167f3ebe[14]),
    .b(al_a352434c[11]),
    .c(al_f57392c),
    .o(al_7452903f[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d63c16e (
    .a(al_167f3ebe[15]),
    .b(al_a352434c[12]),
    .c(al_f57392c),
    .o(al_7452903f[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_615e51b9 (
    .a(al_167f3ebe[16]),
    .b(al_a352434c[13]),
    .c(al_f57392c),
    .o(al_7452903f[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_50f1e904 (
    .a(al_167f3ebe[17]),
    .b(al_a352434c[14]),
    .c(al_f57392c),
    .o(al_7452903f[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_be995e49 (
    .a(al_167f3ebe[18]),
    .b(al_a352434c[15]),
    .c(al_f57392c),
    .o(al_7452903f[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d534c0ef (
    .a(al_167f3ebe[19]),
    .b(al_a352434c[16]),
    .c(al_f57392c),
    .o(al_7452903f[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a3c54db0 (
    .a(al_167f3ebe[20]),
    .b(al_a352434c[17]),
    .c(al_f57392c),
    .o(al_7452903f[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4aef6df3 (
    .a(al_167f3ebe[21]),
    .b(al_a352434c[18]),
    .c(al_f57392c),
    .o(al_7452903f[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_97a2ef97 (
    .a(al_167f3ebe[22]),
    .b(al_a352434c[19]),
    .c(al_f57392c),
    .o(al_7452903f[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_8b9b10e9 (
    .a(al_167f3ebe[23]),
    .b(al_a352434c[20]),
    .c(al_f57392c),
    .o(al_7452903f[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_eb192829 (
    .a(al_167f3ebe[24]),
    .b(al_a352434c[21]),
    .c(al_f57392c),
    .o(al_7452903f[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d97ec514 (
    .a(al_167f3ebe[25]),
    .b(al_a352434c[22]),
    .c(al_f57392c),
    .o(al_7452903f[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5842e8ee (
    .a(al_167f3ebe[26]),
    .b(al_a352434c[23]),
    .c(al_f57392c),
    .o(al_7452903f[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_61e67816 (
    .a(al_167f3ebe[27]),
    .b(al_a352434c[24]),
    .c(al_f57392c),
    .o(al_7452903f[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d3c9b660 (
    .a(al_167f3ebe[28]),
    .b(al_a352434c[25]),
    .c(al_f57392c),
    .o(al_7452903f[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2ee5805a (
    .a(al_167f3ebe[29]),
    .b(al_a352434c[26]),
    .c(al_f57392c),
    .o(al_7452903f[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b3b18589 (
    .a(al_167f3ebe[30]),
    .b(al_a352434c[27]),
    .c(al_f57392c),
    .o(al_7452903f[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9cc001da (
    .a(al_167f3ebe[31]),
    .b(al_a352434c[28]),
    .c(al_f57392c),
    .o(al_7452903f[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1c277e0c (
    .a(al_167f3ebe[32]),
    .b(al_a352434c[29]),
    .c(al_f57392c),
    .o(al_7452903f[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2c261333 (
    .a(al_167f3ebe[33]),
    .b(al_a352434c[30]),
    .c(al_f57392c),
    .o(al_7452903f[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f2ae98d2 (
    .a(al_167f3ebe[34]),
    .b(al_a352434c[31]),
    .c(al_f57392c),
    .o(al_7452903f[34]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_456b48d4 (
    .a(al_167f3ebe[3]),
    .b(al_a352434c[0]),
    .c(al_f57392c),
    .o(al_7452903f[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f49b38ac (
    .a(al_167f3ebe[4]),
    .b(al_a352434c[1]),
    .c(al_f57392c),
    .o(al_7452903f[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d822e846 (
    .a(al_167f3ebe[5]),
    .b(al_a352434c[2]),
    .c(al_f57392c),
    .o(al_7452903f[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4f67acf0 (
    .a(al_167f3ebe[6]),
    .b(al_a352434c[3]),
    .c(al_f57392c),
    .o(al_7452903f[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ff7f5ef9 (
    .a(al_167f3ebe[7]),
    .b(al_a352434c[4]),
    .c(al_f57392c),
    .o(al_7452903f[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_22b8f46d (
    .a(al_167f3ebe[8]),
    .b(al_a352434c[5]),
    .c(al_f57392c),
    .o(al_7452903f[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f8789577 (
    .a(al_167f3ebe[9]),
    .b(al_a352434c[6]),
    .c(al_f57392c),
    .o(al_7452903f[9]));
  AL_DFF_X al_f211b052 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_167f3ebe[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[0]));
  AL_DFF_X al_ab861d64 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[9]));
  AL_DFF_X al_17b0d3b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[10]));
  AL_DFF_X al_b87ff500 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[11]));
  AL_DFF_X al_846ce372 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[12]));
  AL_DFF_X al_e9f517ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[13]));
  AL_DFF_X al_6e17388a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[14]));
  AL_DFF_X al_2ecbe677 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[15]));
  AL_DFF_X al_6070f382 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[16]));
  AL_DFF_X al_918fa82d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[17]));
  AL_DFF_X al_b138f985 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[18]));
  AL_DFF_X al_a5d74aec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_167f3ebe[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[1]));
  AL_DFF_X al_e011a27d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[19]));
  AL_DFF_X al_452d462a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[20]));
  AL_DFF_X al_b06ce9df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[21]));
  AL_DFF_X al_3a91b1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[22]));
  AL_DFF_X al_a45bee8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[23]));
  AL_DFF_X al_a02620b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[24]));
  AL_DFF_X al_ae40b964 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[25]));
  AL_DFF_X al_2bdae326 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[26]));
  AL_DFF_X al_b72fbba6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[27]));
  AL_DFF_X al_f47fb65b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[28]));
  AL_DFF_X al_1cd58229 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_167f3ebe[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[2]));
  AL_DFF_X al_5c9bb3bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[29]));
  AL_DFF_X al_4752cad1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[30]));
  AL_DFF_X al_c40c6c06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[31]));
  AL_DFF_X al_f0058894 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[32]));
  AL_DFF_X al_949334aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[33]));
  AL_DFF_X al_5b300d39 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[34]));
  AL_DFF_X al_c76a137a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[3]));
  AL_DFF_X al_f1cd4ee3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[4]));
  AL_DFF_X al_8e318c10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[5]));
  AL_DFF_X al_7df0df09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[6]));
  AL_DFF_X al_c4a4c5a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[7]));
  AL_DFF_X al_1b4882ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7452903f[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_cafe0ad[8]));
  AL_DFF_X al_d717e864 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f57392c),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[0]));
  AL_DFF_X al_cb119ad8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[9]));
  AL_DFF_X al_be4d628e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[10]));
  AL_DFF_X al_9086ef50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[11]));
  AL_DFF_X al_1ebde988 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[12]));
  AL_DFF_X al_66bb2a18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[13]));
  AL_DFF_X al_f91e4864 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[14]));
  AL_DFF_X al_fe17deee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[15]));
  AL_DFF_X al_96288237 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[16]));
  AL_DFF_X al_21dc34ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[17]));
  AL_DFF_X al_78352827 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[18]));
  AL_DFF_X al_80d938da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[1]));
  AL_DFF_X al_69263dd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[19]));
  AL_DFF_X al_c7b1482c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[20]));
  AL_DFF_X al_c417b7c4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[21]));
  AL_DFF_X al_e0104349 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[22]));
  AL_DFF_X al_960df33a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[23]));
  AL_DFF_X al_8b87b4a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[24]));
  AL_DFF_X al_e63eb7b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[25]));
  AL_DFF_X al_d16052d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[26]));
  AL_DFF_X al_c3a7aec3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[27]));
  AL_DFF_X al_e97ba29f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[28]));
  AL_DFF_X al_aa0f1944 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[2]));
  AL_DFF_X al_1da7c7c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[29]));
  AL_DFF_X al_9f64b116 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[30]));
  AL_DFF_X al_5922ebe1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[31]));
  AL_DFF_X al_5737bfd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[32]));
  AL_DFF_X al_ea055437 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[33]));
  AL_DFF_X al_3fa35306 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[34]));
  AL_DFF_X al_909f91d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[35]));
  AL_DFF_X al_a8d36f53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[36]));
  AL_DFF_X al_bc9de2ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[37]));
  AL_DFF_X al_37520b63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[38]));
  AL_DFF_X al_4b423d52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[3]));
  AL_DFF_X al_876d3bcb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[39]));
  AL_DFF_X al_372fae38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[40]));
  AL_DFF_X al_4b12699e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[41]));
  AL_DFF_X al_2bd024da (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[42]));
  AL_DFF_X al_ea43186 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[43]));
  AL_DFF_X al_f53d39c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[44]));
  AL_DFF_X al_54f4dcb8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[4]));
  AL_DFF_X al_d6a465d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[5]));
  AL_DFF_X al_715dd1a9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[6]));
  AL_DFF_X al_c33358a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[7]));
  AL_DFF_X al_57376d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c2cdf2f1[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_2c312a8[8]));
  AL_DFF_X al_c60a4916 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5d2b923b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1fd6d456[0]));
  AL_DFF_X al_d62d8f9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[9]));
  AL_DFF_X al_ac6e83e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[10]));
  AL_DFF_X al_b471af68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[11]));
  AL_DFF_X al_c1474ab8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[12]));
  AL_DFF_X al_a3cc7f91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[13]));
  AL_DFF_X al_c4a3dbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[14]));
  AL_DFF_X al_d3e2a892 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[15]));
  AL_DFF_X al_295cbd6b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[16]));
  AL_DFF_X al_4fe16805 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[17]));
  AL_DFF_X al_3bc86918 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[18]));
  AL_DFF_X al_1aacf9cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[1]));
  AL_DFF_X al_78b63cc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[19]));
  AL_DFF_X al_f2a55f60 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[20]));
  AL_DFF_X al_8bbc6310 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[21]));
  AL_DFF_X al_f9f50d01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[22]));
  AL_DFF_X al_3f5f749e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[23]));
  AL_DFF_X al_890f97ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[24]));
  AL_DFF_X al_87059e90 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[25]));
  AL_DFF_X al_ea972e88 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[26]));
  AL_DFF_X al_e318afb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[27]));
  AL_DFF_X al_e637d743 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[28]));
  AL_DFF_X al_357730de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[2]));
  AL_DFF_X al_477120c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[29]));
  AL_DFF_X al_214ee352 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[30]));
  AL_DFF_X al_a6ed1986 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[31]));
  AL_DFF_X al_3aca14ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[32]));
  AL_DFF_X al_b1a8b3fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[3]));
  AL_DFF_X al_3c265034 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[4]));
  AL_DFF_X al_3ca0bb32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[5]));
  AL_DFF_X al_c2e22bfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[6]));
  AL_DFF_X al_eefe5917 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[7]));
  AL_DFF_X al_e45d1fe4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7e0865ed[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8ee40da8[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_2fcdc4eb (
    .a(1'b0),
    .o({al_9dc8cf16,open_n197}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bb0c04ae (
    .a(al_cafe0ad[2]),
    .b(al_7e0865ed[2]),
    .c(al_9dc8cf16),
    .o({al_23f7cf96,al_fc56973[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_41d73c0c (
    .a(al_cafe0ad[3]),
    .b(al_7e0865ed[3]),
    .c(al_23f7cf96),
    .o({al_6007eb01,al_fc56973[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dfe59cf0 (
    .a(al_cafe0ad[4]),
    .b(al_7e0865ed[4]),
    .c(al_6007eb01),
    .o({al_e9dcbf51,al_fc56973[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a57ef5e4 (
    .a(al_cafe0ad[5]),
    .b(al_7e0865ed[5]),
    .c(al_e9dcbf51),
    .o({al_af282b4e,al_fc56973[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b3030195 (
    .a(al_cafe0ad[6]),
    .b(al_7e0865ed[6]),
    .c(al_af282b4e),
    .o({al_f13375bf,al_fc56973[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a1a2a809 (
    .a(al_cafe0ad[7]),
    .b(al_7e0865ed[7]),
    .c(al_f13375bf),
    .o({al_79e6f53f,al_fc56973[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_36914fbf (
    .a(al_cafe0ad[8]),
    .b(al_7e0865ed[8]),
    .c(al_79e6f53f),
    .o({al_262f4fd9,al_fc56973[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_de03aaea (
    .a(al_cafe0ad[9]),
    .b(al_7e0865ed[9]),
    .c(al_262f4fd9),
    .o({al_91a1715,al_fc56973[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6f7e7ed0 (
    .a(al_cafe0ad[10]),
    .b(al_7e0865ed[10]),
    .c(al_91a1715),
    .o({al_466678a0,al_fc56973[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3825ac92 (
    .a(al_cafe0ad[11]),
    .b(al_7e0865ed[11]),
    .c(al_466678a0),
    .o({al_b3412438,al_fc56973[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8ddb8883 (
    .a(al_cafe0ad[12]),
    .b(al_7e0865ed[12]),
    .c(al_b3412438),
    .o({al_905abb5d,al_fc56973[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c0ceb33b (
    .a(al_cafe0ad[13]),
    .b(al_7e0865ed[13]),
    .c(al_905abb5d),
    .o({al_30d2d597,al_fc56973[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f17f3fab (
    .a(al_cafe0ad[14]),
    .b(al_7e0865ed[14]),
    .c(al_30d2d597),
    .o({al_b4ebcfb5,al_fc56973[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7dc6aa19 (
    .a(al_cafe0ad[15]),
    .b(al_7e0865ed[15]),
    .c(al_b4ebcfb5),
    .o({al_9398f98d,al_fc56973[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6bd4991d (
    .a(al_cafe0ad[16]),
    .b(al_7e0865ed[16]),
    .c(al_9398f98d),
    .o({al_2e77c07b,al_fc56973[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c2d78f9b (
    .a(al_cafe0ad[17]),
    .b(al_7e0865ed[17]),
    .c(al_2e77c07b),
    .o({al_56c765b9,al_fc56973[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b30ca66e (
    .a(al_cafe0ad[18]),
    .b(al_7e0865ed[18]),
    .c(al_56c765b9),
    .o({al_abeeae47,al_fc56973[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_61e495a7 (
    .a(al_cafe0ad[19]),
    .b(al_7e0865ed[19]),
    .c(al_abeeae47),
    .o({al_59c21146,al_fc56973[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1fee88dc (
    .a(al_cafe0ad[20]),
    .b(al_7e0865ed[20]),
    .c(al_59c21146),
    .o({al_e154cc8,al_fc56973[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a690a852 (
    .a(al_cafe0ad[21]),
    .b(al_7e0865ed[21]),
    .c(al_e154cc8),
    .o({al_c2370696,al_fc56973[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2a5af59a (
    .a(al_cafe0ad[22]),
    .b(al_7e0865ed[22]),
    .c(al_c2370696),
    .o({al_c0c45a44,al_fc56973[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_37bc3c3c (
    .a(al_cafe0ad[23]),
    .b(al_7e0865ed[23]),
    .c(al_c0c45a44),
    .o({al_32d5e65b,al_fc56973[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_83f5558a (
    .a(al_cafe0ad[24]),
    .b(al_7e0865ed[24]),
    .c(al_32d5e65b),
    .o({al_627e2733,al_fc56973[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c931e3ed (
    .a(al_cafe0ad[25]),
    .b(al_7e0865ed[25]),
    .c(al_627e2733),
    .o({al_4caf87a4,al_fc56973[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4882656 (
    .a(al_cafe0ad[26]),
    .b(al_7e0865ed[26]),
    .c(al_4caf87a4),
    .o({al_93eba83e,al_fc56973[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_85ca9881 (
    .a(al_cafe0ad[27]),
    .b(al_7e0865ed[27]),
    .c(al_93eba83e),
    .o({al_f4b95543,al_fc56973[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2c04c1b7 (
    .a(al_cafe0ad[28]),
    .b(al_7e0865ed[28]),
    .c(al_f4b95543),
    .o({al_431d20ff,al_fc56973[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ec0e437c (
    .a(al_cafe0ad[29]),
    .b(al_7e0865ed[29]),
    .c(al_431d20ff),
    .o({al_12da8cbc,al_fc56973[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9b46f2c6 (
    .a(al_cafe0ad[30]),
    .b(al_7e0865ed[30]),
    .c(al_12da8cbc),
    .o({al_a05b5ad4,al_fc56973[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b81de1e7 (
    .a(al_cafe0ad[31]),
    .b(al_7e0865ed[31]),
    .c(al_a05b5ad4),
    .o({al_5072fc21,al_fc56973[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_92554506 (
    .a(al_cafe0ad[32]),
    .b(al_7e0865ed[32]),
    .c(al_5072fc21),
    .o({al_e6b19e19,al_fc56973[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e0cfd00a (
    .a(al_cafe0ad[33]),
    .b(al_7e0865ed[33]),
    .c(al_e6b19e19),
    .o({al_baadae4d,al_fc56973[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1bf1c0b8 (
    .a(al_cafe0ad[34]),
    .b(1'b0),
    .c(al_baadae4d),
    .o({al_c4be0e1d,open_n198}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_754c2ef8 (
    .a(1'b0),
    .b(1'b1),
    .c(al_c4be0e1d),
    .o({open_n199,al_5dc8be80}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_2faa16fe (
    .a(al_cafe0ad[10]),
    .b(al_fc56973[8]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_68a2008c (
    .a(al_cafe0ad[11]),
    .b(al_fc56973[9]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bad8f580 (
    .a(al_cafe0ad[12]),
    .b(al_fc56973[10]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5b798a6 (
    .a(al_cafe0ad[13]),
    .b(al_fc56973[11]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3be796f7 (
    .a(al_cafe0ad[14]),
    .b(al_fc56973[12]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ad859397 (
    .a(al_cafe0ad[15]),
    .b(al_fc56973[13]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_98fb5936 (
    .a(al_cafe0ad[16]),
    .b(al_fc56973[14]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7b967c60 (
    .a(al_cafe0ad[17]),
    .b(al_fc56973[15]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_42ed5e3c (
    .a(al_cafe0ad[18]),
    .b(al_fc56973[16]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cbd5c5c2 (
    .a(al_cafe0ad[19]),
    .b(al_fc56973[17]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bf52eee9 (
    .a(al_cafe0ad[20]),
    .b(al_fc56973[18]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f49edfa8 (
    .a(al_cafe0ad[21]),
    .b(al_fc56973[19]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_caced78 (
    .a(al_cafe0ad[22]),
    .b(al_fc56973[20]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_54205bdb (
    .a(al_cafe0ad[23]),
    .b(al_fc56973[21]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3163d62d (
    .a(al_cafe0ad[24]),
    .b(al_fc56973[22]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a14deecd (
    .a(al_cafe0ad[25]),
    .b(al_fc56973[23]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3328429f (
    .a(al_cafe0ad[26]),
    .b(al_fc56973[24]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1e28ec86 (
    .a(al_cafe0ad[27]),
    .b(al_fc56973[25]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_92e03d9 (
    .a(al_cafe0ad[28]),
    .b(al_fc56973[26]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b1a7dba5 (
    .a(al_cafe0ad[29]),
    .b(al_fc56973[27]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_74fa56a3 (
    .a(al_cafe0ad[2]),
    .b(al_fc56973[0]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d310dff (
    .a(al_cafe0ad[30]),
    .b(al_fc56973[28]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_edf77648 (
    .a(al_cafe0ad[31]),
    .b(al_fc56973[29]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e9815af0 (
    .a(al_cafe0ad[32]),
    .b(al_fc56973[30]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f66d6bc1 (
    .a(al_cafe0ad[33]),
    .b(al_fc56973[31]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[33]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9417d59c (
    .a(al_cafe0ad[3]),
    .b(al_fc56973[1]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f45823ff (
    .a(al_cafe0ad[4]),
    .b(al_fc56973[2]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_39fc5f85 (
    .a(al_cafe0ad[5]),
    .b(al_fc56973[3]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e77967d1 (
    .a(al_cafe0ad[6]),
    .b(al_fc56973[4]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_817f5204 (
    .a(al_cafe0ad[7]),
    .b(al_fc56973[5]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_25c3dedc (
    .a(al_cafe0ad[8]),
    .b(al_fc56973[6]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_577b734a (
    .a(al_cafe0ad[9]),
    .b(al_fc56973[7]),
    .c(al_5dc8be80),
    .o(al_ce2f96cc[9]));
  AL_DFF_X al_e33da38 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cafe0ad[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[0]));
  AL_DFF_X al_76d79639 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[9]));
  AL_DFF_X al_871e1cc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[10]));
  AL_DFF_X al_98e7d3ed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[11]));
  AL_DFF_X al_ea64b014 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[12]));
  AL_DFF_X al_1e74ef43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[13]));
  AL_DFF_X al_db832f3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[14]));
  AL_DFF_X al_a1f3ec02 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[15]));
  AL_DFF_X al_403b3694 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[16]));
  AL_DFF_X al_fbdb3203 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[17]));
  AL_DFF_X al_7cfad07 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[18]));
  AL_DFF_X al_ddeb37a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_cafe0ad[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[1]));
  AL_DFF_X al_eb993414 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[19]));
  AL_DFF_X al_b071220c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[20]));
  AL_DFF_X al_7eaa75b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[21]));
  AL_DFF_X al_a7ed1218 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[22]));
  AL_DFF_X al_d7dfe5b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[23]));
  AL_DFF_X al_665b8b87 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[24]));
  AL_DFF_X al_abc38db4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[25]));
  AL_DFF_X al_5acbb98b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[26]));
  AL_DFF_X al_b3c619e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[27]));
  AL_DFF_X al_d525a8be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[28]));
  AL_DFF_X al_d4160540 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[2]));
  AL_DFF_X al_b14b3cef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[29]));
  AL_DFF_X al_68b4e327 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[30]));
  AL_DFF_X al_aa171412 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[31]));
  AL_DFF_X al_818c2872 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[32]));
  AL_DFF_X al_e7c97f7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[33]));
  AL_DFF_X al_af9d4d48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[3]));
  AL_DFF_X al_2456c61a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[4]));
  AL_DFF_X al_f4384747 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[5]));
  AL_DFF_X al_cd8829ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[6]));
  AL_DFF_X al_aa4d8cbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[7]));
  AL_DFF_X al_b31aa445 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_ce2f96cc[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_13d036ce[8]));
  AL_DFF_X al_5fa73810 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5dc8be80),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[0]));
  AL_DFF_X al_7b992167 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[9]));
  AL_DFF_X al_ec0de4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[10]));
  AL_DFF_X al_48bb09c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[11]));
  AL_DFF_X al_736752fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[12]));
  AL_DFF_X al_768951bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[13]));
  AL_DFF_X al_b806116d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[14]));
  AL_DFF_X al_289cddae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[15]));
  AL_DFF_X al_4888f166 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[16]));
  AL_DFF_X al_a959883f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[17]));
  AL_DFF_X al_1ffd0add (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[18]));
  AL_DFF_X al_7c2e5920 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[1]));
  AL_DFF_X al_8de780c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[19]));
  AL_DFF_X al_1483c033 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[20]));
  AL_DFF_X al_cfb10b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[21]));
  AL_DFF_X al_614f4a54 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[22]));
  AL_DFF_X al_3ce64e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[23]));
  AL_DFF_X al_7fca690c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[24]));
  AL_DFF_X al_6ce0df79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[25]));
  AL_DFF_X al_cb947976 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[26]));
  AL_DFF_X al_f84c4c7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[27]));
  AL_DFF_X al_a4b94f1e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[28]));
  AL_DFF_X al_9730ec0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[2]));
  AL_DFF_X al_cc00df0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[29]));
  AL_DFF_X al_d4039180 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[30]));
  AL_DFF_X al_f5111680 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[31]));
  AL_DFF_X al_828cd183 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[32]));
  AL_DFF_X al_28c846e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[33]));
  AL_DFF_X al_d3f75ccf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[34]));
  AL_DFF_X al_7a79eda9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[35]));
  AL_DFF_X al_a466f790 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[36]));
  AL_DFF_X al_337d25ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[37]));
  AL_DFF_X al_94050b9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[38]));
  AL_DFF_X al_fd32ab16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[3]));
  AL_DFF_X al_1e1f5565 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[39]));
  AL_DFF_X al_3aca2f53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[40]));
  AL_DFF_X al_3abb4cd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[41]));
  AL_DFF_X al_ad51fa31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[42]));
  AL_DFF_X al_f8f37573 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[43]));
  AL_DFF_X al_2d573722 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[44]));
  AL_DFF_X al_c5719f79 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[45]));
  AL_DFF_X al_6b621b72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[4]));
  AL_DFF_X al_c7734ad1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[5]));
  AL_DFF_X al_d5375b91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[6]));
  AL_DFF_X al_3abfec58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[7]));
  AL_DFF_X al_a4a84820 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_2c312a8[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f3197cbe[8]));
  AL_DFF_X al_994632cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1fd6d456[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_7a934789[0]));
  AL_DFF_X al_b4687cf6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[0]));
  AL_DFF_X al_812802a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[9]));
  AL_DFF_X al_75a98e51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[10]));
  AL_DFF_X al_69622cd5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[11]));
  AL_DFF_X al_53cf3e19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[12]));
  AL_DFF_X al_90175a16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[13]));
  AL_DFF_X al_f74b3c51 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[14]));
  AL_DFF_X al_d735990a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[15]));
  AL_DFF_X al_aa8175eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[16]));
  AL_DFF_X al_12cec144 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[17]));
  AL_DFF_X al_3026e6e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[18]));
  AL_DFF_X al_ef9bdae2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[1]));
  AL_DFF_X al_274b3bb5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[19]));
  AL_DFF_X al_356d9c41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[20]));
  AL_DFF_X al_946f4700 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[21]));
  AL_DFF_X al_19958099 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[22]));
  AL_DFF_X al_767651e3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[23]));
  AL_DFF_X al_778bb58e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[24]));
  AL_DFF_X al_3d92daee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[25]));
  AL_DFF_X al_4f8eee63 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[26]));
  AL_DFF_X al_f39e296d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[27]));
  AL_DFF_X al_6cc92aef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[28]));
  AL_DFF_X al_24d3ea33 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[2]));
  AL_DFF_X al_34eca8d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[29]));
  AL_DFF_X al_817f4dbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[30]));
  AL_DFF_X al_23dee699 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[31]));
  AL_DFF_X al_4a17483c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[3]));
  AL_DFF_X al_9780161e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[4]));
  AL_DFF_X al_5e74f527 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[5]));
  AL_DFF_X al_ea67f81b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[6]));
  AL_DFF_X al_f87896de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[7]));
  AL_DFF_X al_42b1d803 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8ee40da8[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_ac1cba4d[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_6595569e (
    .a(1'b0),
    .o({al_547ff558,open_n202}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8dc78814 (
    .a(al_13d036ce[1]),
    .b(al_8ee40da8[1]),
    .c(al_547ff558),
    .o({al_ecd1dd20,al_65caf2b5[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_475a140b (
    .a(al_13d036ce[2]),
    .b(al_8ee40da8[2]),
    .c(al_ecd1dd20),
    .o({al_a4a9db62,al_65caf2b5[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27a39a3a (
    .a(al_13d036ce[3]),
    .b(al_8ee40da8[3]),
    .c(al_a4a9db62),
    .o({al_2150e0ab,al_65caf2b5[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b8a2a191 (
    .a(al_13d036ce[4]),
    .b(al_8ee40da8[4]),
    .c(al_2150e0ab),
    .o({al_98763df0,al_65caf2b5[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f3f482a6 (
    .a(al_13d036ce[5]),
    .b(al_8ee40da8[5]),
    .c(al_98763df0),
    .o({al_a2aa2d49,al_65caf2b5[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_80ded82c (
    .a(al_13d036ce[6]),
    .b(al_8ee40da8[6]),
    .c(al_a2aa2d49),
    .o({al_e749a18b,al_65caf2b5[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e7a9ff08 (
    .a(al_13d036ce[7]),
    .b(al_8ee40da8[7]),
    .c(al_e749a18b),
    .o({al_65250a4c,al_65caf2b5[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_74db9c85 (
    .a(al_13d036ce[8]),
    .b(al_8ee40da8[8]),
    .c(al_65250a4c),
    .o({al_71dba21f,al_65caf2b5[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_6208bf58 (
    .a(al_13d036ce[9]),
    .b(al_8ee40da8[9]),
    .c(al_71dba21f),
    .o({al_5ba1798e,al_65caf2b5[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1c0583ff (
    .a(al_13d036ce[10]),
    .b(al_8ee40da8[10]),
    .c(al_5ba1798e),
    .o({al_fa3cfc2c,al_65caf2b5[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ea13415e (
    .a(al_13d036ce[11]),
    .b(al_8ee40da8[11]),
    .c(al_fa3cfc2c),
    .o({al_eebdc4f4,al_65caf2b5[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b009c1d1 (
    .a(al_13d036ce[12]),
    .b(al_8ee40da8[12]),
    .c(al_eebdc4f4),
    .o({al_88900ac6,al_65caf2b5[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ddcdc003 (
    .a(al_13d036ce[13]),
    .b(al_8ee40da8[13]),
    .c(al_88900ac6),
    .o({al_f1ea9238,al_65caf2b5[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ef527df7 (
    .a(al_13d036ce[14]),
    .b(al_8ee40da8[14]),
    .c(al_f1ea9238),
    .o({al_cb718520,al_65caf2b5[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_425124d3 (
    .a(al_13d036ce[15]),
    .b(al_8ee40da8[15]),
    .c(al_cb718520),
    .o({al_47b988e0,al_65caf2b5[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c2116d73 (
    .a(al_13d036ce[16]),
    .b(al_8ee40da8[16]),
    .c(al_47b988e0),
    .o({al_919eb56e,al_65caf2b5[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_322e6a6c (
    .a(al_13d036ce[17]),
    .b(al_8ee40da8[17]),
    .c(al_919eb56e),
    .o({al_35e6fce8,al_65caf2b5[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e583fa8e (
    .a(al_13d036ce[18]),
    .b(al_8ee40da8[18]),
    .c(al_35e6fce8),
    .o({al_6a0855b2,al_65caf2b5[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c6c26b9b (
    .a(al_13d036ce[19]),
    .b(al_8ee40da8[19]),
    .c(al_6a0855b2),
    .o({al_607eee13,al_65caf2b5[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bdef8cf1 (
    .a(al_13d036ce[20]),
    .b(al_8ee40da8[20]),
    .c(al_607eee13),
    .o({al_9f13bda9,al_65caf2b5[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b494ad9 (
    .a(al_13d036ce[21]),
    .b(al_8ee40da8[21]),
    .c(al_9f13bda9),
    .o({al_7d943beb,al_65caf2b5[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9c407d0b (
    .a(al_13d036ce[22]),
    .b(al_8ee40da8[22]),
    .c(al_7d943beb),
    .o({al_6d747586,al_65caf2b5[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_264d183d (
    .a(al_13d036ce[23]),
    .b(al_8ee40da8[23]),
    .c(al_6d747586),
    .o({al_d6a2647c,al_65caf2b5[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc9bc59c (
    .a(al_13d036ce[24]),
    .b(al_8ee40da8[24]),
    .c(al_d6a2647c),
    .o({al_8cb59e89,al_65caf2b5[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3fa06b6b (
    .a(al_13d036ce[25]),
    .b(al_8ee40da8[25]),
    .c(al_8cb59e89),
    .o({al_63e85dd3,al_65caf2b5[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2c640d7 (
    .a(al_13d036ce[26]),
    .b(al_8ee40da8[26]),
    .c(al_63e85dd3),
    .o({al_2d304c84,al_65caf2b5[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c9e1f963 (
    .a(al_13d036ce[27]),
    .b(al_8ee40da8[27]),
    .c(al_2d304c84),
    .o({al_59db63b2,al_65caf2b5[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3dde0dc2 (
    .a(al_13d036ce[28]),
    .b(al_8ee40da8[28]),
    .c(al_59db63b2),
    .o({al_ef9e6ec2,al_65caf2b5[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8d6ed8db (
    .a(al_13d036ce[29]),
    .b(al_8ee40da8[29]),
    .c(al_ef9e6ec2),
    .o({al_ee134d8c,al_65caf2b5[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3f2c1c9b (
    .a(al_13d036ce[30]),
    .b(al_8ee40da8[30]),
    .c(al_ee134d8c),
    .o({al_931bfadf,al_65caf2b5[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_40467f7e (
    .a(al_13d036ce[31]),
    .b(al_8ee40da8[31]),
    .c(al_931bfadf),
    .o({al_f57240df,al_65caf2b5[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b1577177 (
    .a(al_13d036ce[32]),
    .b(al_8ee40da8[32]),
    .c(al_f57240df),
    .o({al_d1cf7fc7,al_65caf2b5[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_16c8b487 (
    .a(al_13d036ce[33]),
    .b(1'b0),
    .c(al_d1cf7fc7),
    .o({al_f80ea3fa,open_n203}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_27b5bc17 (
    .a(1'b0),
    .b(1'b1),
    .c(al_f80ea3fa),
    .o({open_n204,al_6cebde96}));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6dd95848 (
    .a(al_13d036ce[10]),
    .b(al_65caf2b5[9]),
    .c(al_6cebde96),
    .o(al_b328a515[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f63966ab (
    .a(al_13d036ce[11]),
    .b(al_65caf2b5[10]),
    .c(al_6cebde96),
    .o(al_b328a515[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_21bc7845 (
    .a(al_13d036ce[12]),
    .b(al_65caf2b5[11]),
    .c(al_6cebde96),
    .o(al_b328a515[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ea4fc59e (
    .a(al_13d036ce[13]),
    .b(al_65caf2b5[12]),
    .c(al_6cebde96),
    .o(al_b328a515[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_97456e0 (
    .a(al_13d036ce[14]),
    .b(al_65caf2b5[13]),
    .c(al_6cebde96),
    .o(al_b328a515[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_4bf4072e (
    .a(al_13d036ce[15]),
    .b(al_65caf2b5[14]),
    .c(al_6cebde96),
    .o(al_b328a515[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9c33f903 (
    .a(al_13d036ce[16]),
    .b(al_65caf2b5[15]),
    .c(al_6cebde96),
    .o(al_b328a515[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fbf52dd0 (
    .a(al_13d036ce[17]),
    .b(al_65caf2b5[16]),
    .c(al_6cebde96),
    .o(al_b328a515[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ce4d7c5f (
    .a(al_13d036ce[18]),
    .b(al_65caf2b5[17]),
    .c(al_6cebde96),
    .o(al_b328a515[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f8585708 (
    .a(al_13d036ce[19]),
    .b(al_65caf2b5[18]),
    .c(al_6cebde96),
    .o(al_b328a515[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_bf1a6718 (
    .a(al_13d036ce[1]),
    .b(al_65caf2b5[0]),
    .c(al_6cebde96),
    .o(al_b328a515[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a7bc501d (
    .a(al_13d036ce[20]),
    .b(al_65caf2b5[19]),
    .c(al_6cebde96),
    .o(al_b328a515[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a519e0bd (
    .a(al_13d036ce[21]),
    .b(al_65caf2b5[20]),
    .c(al_6cebde96),
    .o(al_b328a515[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3f79db9c (
    .a(al_13d036ce[22]),
    .b(al_65caf2b5[21]),
    .c(al_6cebde96),
    .o(al_b328a515[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_9965cf06 (
    .a(al_13d036ce[23]),
    .b(al_65caf2b5[22]),
    .c(al_6cebde96),
    .o(al_b328a515[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3bddf734 (
    .a(al_13d036ce[24]),
    .b(al_65caf2b5[23]),
    .c(al_6cebde96),
    .o(al_b328a515[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5f2e0e3 (
    .a(al_13d036ce[25]),
    .b(al_65caf2b5[24]),
    .c(al_6cebde96),
    .o(al_b328a515[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e5b88769 (
    .a(al_13d036ce[26]),
    .b(al_65caf2b5[25]),
    .c(al_6cebde96),
    .o(al_b328a515[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5b3666d1 (
    .a(al_13d036ce[27]),
    .b(al_65caf2b5[26]),
    .c(al_6cebde96),
    .o(al_b328a515[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_af9271c (
    .a(al_13d036ce[28]),
    .b(al_65caf2b5[27]),
    .c(al_6cebde96),
    .o(al_b328a515[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_f95f9197 (
    .a(al_13d036ce[29]),
    .b(al_65caf2b5[28]),
    .c(al_6cebde96),
    .o(al_b328a515[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6a250738 (
    .a(al_13d036ce[2]),
    .b(al_65caf2b5[1]),
    .c(al_6cebde96),
    .o(al_b328a515[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ca063cef (
    .a(al_13d036ce[30]),
    .b(al_65caf2b5[29]),
    .c(al_6cebde96),
    .o(al_b328a515[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6af2d1da (
    .a(al_13d036ce[31]),
    .b(al_65caf2b5[30]),
    .c(al_6cebde96),
    .o(al_b328a515[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b84eac01 (
    .a(al_13d036ce[32]),
    .b(al_65caf2b5[31]),
    .c(al_6cebde96),
    .o(al_b328a515[32]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_20db0a84 (
    .a(al_13d036ce[3]),
    .b(al_65caf2b5[2]),
    .c(al_6cebde96),
    .o(al_b328a515[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_79314098 (
    .a(al_13d036ce[4]),
    .b(al_65caf2b5[3]),
    .c(al_6cebde96),
    .o(al_b328a515[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a7770fdf (
    .a(al_13d036ce[5]),
    .b(al_65caf2b5[4]),
    .c(al_6cebde96),
    .o(al_b328a515[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3779d4be (
    .a(al_13d036ce[6]),
    .b(al_65caf2b5[5]),
    .c(al_6cebde96),
    .o(al_b328a515[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_30a31136 (
    .a(al_13d036ce[7]),
    .b(al_65caf2b5[6]),
    .c(al_6cebde96),
    .o(al_b328a515[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c6625f89 (
    .a(al_13d036ce[8]),
    .b(al_65caf2b5[7]),
    .c(al_6cebde96),
    .o(al_b328a515[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a4655937 (
    .a(al_13d036ce[9]),
    .b(al_65caf2b5[8]),
    .c(al_6cebde96),
    .o(al_b328a515[9]));
  AL_DFF_X al_980b2d44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_13d036ce[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[0]));
  AL_DFF_X al_89a0398f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[9]));
  AL_DFF_X al_9486c8fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[10]));
  AL_DFF_X al_6e2819db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[11]));
  AL_DFF_X al_a6b6a067 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[12]));
  AL_DFF_X al_56369cac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[13]));
  AL_DFF_X al_17439215 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[14]));
  AL_DFF_X al_514ba8ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[15]));
  AL_DFF_X al_d2ccda5f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[16]));
  AL_DFF_X al_f433a28f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[17]));
  AL_DFF_X al_3d434ec9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[18]));
  AL_DFF_X al_28c1e1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[1]));
  AL_DFF_X al_91e5405c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[19]));
  AL_DFF_X al_67944697 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[20]));
  AL_DFF_X al_bb9928d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[21]));
  AL_DFF_X al_b5a05793 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[22]));
  AL_DFF_X al_f8489915 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[23]));
  AL_DFF_X al_d2da9295 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[24]));
  AL_DFF_X al_b31aad58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[25]));
  AL_DFF_X al_3f874cc5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[26]));
  AL_DFF_X al_e9f55e8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[27]));
  AL_DFF_X al_4ae80715 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[28]));
  AL_DFF_X al_6c252d8b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[2]));
  AL_DFF_X al_188d5c1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[29]));
  AL_DFF_X al_2fbfe5f8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[30]));
  AL_DFF_X al_62acb3b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[31]));
  AL_DFF_X al_c49759bd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[32]));
  AL_DFF_X al_ff4678b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[3]));
  AL_DFF_X al_2445a6c3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[4]));
  AL_DFF_X al_47e92470 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[5]));
  AL_DFF_X al_e85fe617 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[6]));
  AL_DFF_X al_39fb17ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[7]));
  AL_DFF_X al_e19979bc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b328a515[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_8f041238[8]));
  AL_DFF_X al_f97a6f15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6cebde96),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[0]));
  AL_DFF_X al_fb5653ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[9]));
  AL_DFF_X al_2692b857 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[10]));
  AL_DFF_X al_8dd1d328 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[11]));
  AL_DFF_X al_ccb52d1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[12]));
  AL_DFF_X al_2e8925f9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[13]));
  AL_DFF_X al_1e1cb986 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[14]));
  AL_DFF_X al_f767c7df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[15]));
  AL_DFF_X al_6339daa0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[16]));
  AL_DFF_X al_817e0b78 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[17]));
  AL_DFF_X al_e2c7f984 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[18]));
  AL_DFF_X al_35ec32a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[1]));
  AL_DFF_X al_4d459a99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[19]));
  AL_DFF_X al_8044581d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[20]));
  AL_DFF_X al_2f4c33d4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[21]));
  AL_DFF_X al_d0403799 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[22]));
  AL_DFF_X al_e04df6f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[23]));
  AL_DFF_X al_b124c91b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[24]));
  AL_DFF_X al_bb6fedfb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[25]));
  AL_DFF_X al_d596e649 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[26]));
  AL_DFF_X al_191e42e5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[27]));
  AL_DFF_X al_5a263280 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[28]));
  AL_DFF_X al_c2b7b3be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[2]));
  AL_DFF_X al_2c618e7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[29]));
  AL_DFF_X al_ec67d055 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[30]));
  AL_DFF_X al_13eb601a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[31]));
  AL_DFF_X al_315c832f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[32]));
  AL_DFF_X al_4bb9c1cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[33]));
  AL_DFF_X al_b7f5ab7d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[34]));
  AL_DFF_X al_c7b63e3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[35]));
  AL_DFF_X al_65086e6c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[36]));
  AL_DFF_X al_8a72b6a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[37]));
  AL_DFF_X al_c3ca7f17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[38]));
  AL_DFF_X al_bab29c1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[3]));
  AL_DFF_X al_2cad2154 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[39]));
  AL_DFF_X al_c87cdb2d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[40]));
  AL_DFF_X al_4c8dd47c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[41]));
  AL_DFF_X al_db622ef7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[42]));
  AL_DFF_X al_4b997766 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[43]));
  AL_DFF_X al_c5e0615 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[44]));
  AL_DFF_X al_5988a191 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[45]));
  AL_DFF_X al_ba5b106 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[46]));
  AL_DFF_X al_1e7d6f70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[4]));
  AL_DFF_X al_78d372c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[5]));
  AL_DFF_X al_4f93f2bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[6]));
  AL_DFF_X al_5c58b4aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[7]));
  AL_DFF_X al_b81907ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f3197cbe[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59124752[8]));
  AL_DFF_X al_955c37fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a934789[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_dc871c53[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e538579b (
    .a(al_8f041238[0]),
    .b(al_42247ac7[0]),
    .c(al_b84db2a6),
    .o(al_4101ed12[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_7b47fb2b (
    .a(al_8f041238[10]),
    .b(al_42247ac7[10]),
    .c(al_b84db2a6),
    .o(al_4101ed12[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_58ffa7f5 (
    .a(al_8f041238[11]),
    .b(al_42247ac7[11]),
    .c(al_b84db2a6),
    .o(al_4101ed12[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c9f4842d (
    .a(al_8f041238[12]),
    .b(al_42247ac7[12]),
    .c(al_b84db2a6),
    .o(al_4101ed12[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_20eb671d (
    .a(al_8f041238[13]),
    .b(al_42247ac7[13]),
    .c(al_b84db2a6),
    .o(al_4101ed12[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_b43001df (
    .a(al_8f041238[14]),
    .b(al_42247ac7[14]),
    .c(al_b84db2a6),
    .o(al_4101ed12[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_20c2bc95 (
    .a(al_8f041238[15]),
    .b(al_42247ac7[15]),
    .c(al_b84db2a6),
    .o(al_4101ed12[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_cd69bd4 (
    .a(al_8f041238[16]),
    .b(al_42247ac7[16]),
    .c(al_b84db2a6),
    .o(al_4101ed12[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_5aeb1b6c (
    .a(al_8f041238[17]),
    .b(al_42247ac7[17]),
    .c(al_b84db2a6),
    .o(al_4101ed12[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_865b209 (
    .a(al_8f041238[18]),
    .b(al_42247ac7[18]),
    .c(al_b84db2a6),
    .o(al_4101ed12[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_1ec43e90 (
    .a(al_8f041238[19]),
    .b(al_42247ac7[19]),
    .c(al_b84db2a6),
    .o(al_4101ed12[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ec6cbd9f (
    .a(al_8f041238[1]),
    .b(al_42247ac7[1]),
    .c(al_b84db2a6),
    .o(al_4101ed12[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_12fd1217 (
    .a(al_8f041238[20]),
    .b(al_42247ac7[20]),
    .c(al_b84db2a6),
    .o(al_4101ed12[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6b253ea2 (
    .a(al_8f041238[21]),
    .b(al_42247ac7[21]),
    .c(al_b84db2a6),
    .o(al_4101ed12[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a8b4c135 (
    .a(al_8f041238[22]),
    .b(al_42247ac7[22]),
    .c(al_b84db2a6),
    .o(al_4101ed12[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_a9923f48 (
    .a(al_8f041238[23]),
    .b(al_42247ac7[23]),
    .c(al_b84db2a6),
    .o(al_4101ed12[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_182a1553 (
    .a(al_8f041238[24]),
    .b(al_42247ac7[24]),
    .c(al_b84db2a6),
    .o(al_4101ed12[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_6485a24 (
    .a(al_8f041238[25]),
    .b(al_42247ac7[25]),
    .c(al_b84db2a6),
    .o(al_4101ed12[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_84503460 (
    .a(al_8f041238[26]),
    .b(al_42247ac7[26]),
    .c(al_b84db2a6),
    .o(al_4101ed12[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_37b29d59 (
    .a(al_8f041238[27]),
    .b(al_42247ac7[27]),
    .c(al_b84db2a6),
    .o(al_4101ed12[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_583ca1f9 (
    .a(al_8f041238[28]),
    .b(al_42247ac7[28]),
    .c(al_b84db2a6),
    .o(al_4101ed12[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_dfbc37df (
    .a(al_8f041238[29]),
    .b(al_42247ac7[29]),
    .c(al_b84db2a6),
    .o(al_4101ed12[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_c971a95b (
    .a(al_8f041238[2]),
    .b(al_42247ac7[2]),
    .c(al_b84db2a6),
    .o(al_4101ed12[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e38c561b (
    .a(al_8f041238[30]),
    .b(al_42247ac7[30]),
    .c(al_b84db2a6),
    .o(al_4101ed12[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_fde49e17 (
    .a(al_8f041238[31]),
    .b(al_42247ac7[31]),
    .c(al_b84db2a6),
    .o(al_4101ed12[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d5f411fe (
    .a(al_8f041238[3]),
    .b(al_42247ac7[3]),
    .c(al_b84db2a6),
    .o(al_4101ed12[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_e0df35c6 (
    .a(al_8f041238[4]),
    .b(al_42247ac7[4]),
    .c(al_b84db2a6),
    .o(al_4101ed12[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_3fa5bb76 (
    .a(al_8f041238[5]),
    .b(al_42247ac7[5]),
    .c(al_b84db2a6),
    .o(al_4101ed12[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_62b67da9 (
    .a(al_8f041238[6]),
    .b(al_42247ac7[6]),
    .c(al_b84db2a6),
    .o(al_4101ed12[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_ecd62940 (
    .a(al_8f041238[7]),
    .b(al_42247ac7[7]),
    .c(al_b84db2a6),
    .o(al_4101ed12[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_d4387f45 (
    .a(al_8f041238[8]),
    .b(al_42247ac7[8]),
    .c(al_b84db2a6),
    .o(al_4101ed12[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    al_222ffc5c (
    .a(al_8f041238[9]),
    .b(al_42247ac7[9]),
    .c(al_b84db2a6),
    .o(al_4101ed12[9]));
  AL_DFF_X al_2988e194 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[0]));
  AL_DFF_X al_e6a2cba8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[9]));
  AL_DFF_X al_474cc38c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[10]));
  AL_DFF_X al_b08ee0de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[11]));
  AL_DFF_X al_f83dbde8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[12]));
  AL_DFF_X al_e389cc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[13]));
  AL_DFF_X al_1385c202 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[14]));
  AL_DFF_X al_fadf88e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[15]));
  AL_DFF_X al_8719dcb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[16]));
  AL_DFF_X al_5165207f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[17]));
  AL_DFF_X al_a9489e0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[18]));
  AL_DFF_X al_bf8cedec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[1]));
  AL_DFF_X al_f9f2de62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[19]));
  AL_DFF_X al_7e145c4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[20]));
  AL_DFF_X al_22b897f1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[21]));
  AL_DFF_X al_e5d8c3e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[22]));
  AL_DFF_X al_76a2d1a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[23]));
  AL_DFF_X al_ff5f895b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[24]));
  AL_DFF_X al_c76e4b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[25]));
  AL_DFF_X al_4244a5a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[26]));
  AL_DFF_X al_531f3bc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[27]));
  AL_DFF_X al_18d0478b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[28]));
  AL_DFF_X al_a63c968e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[2]));
  AL_DFF_X al_5539666e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[29]));
  AL_DFF_X al_fc2d4d85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[30]));
  AL_DFF_X al_50469946 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[31]));
  AL_DFF_X al_59091459 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[3]));
  AL_DFF_X al_8ac589b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[4]));
  AL_DFF_X al_1c448d27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[5]));
  AL_DFF_X al_da9e225 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[6]));
  AL_DFF_X al_ad98bf7e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[7]));
  AL_DFF_X al_6fafddc6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4101ed12[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_bfaf4e7[8]));
  AL_DFF_X al_10ed571d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b84db2a6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[0]));
  AL_DFF_X al_c5d35c14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[9]));
  AL_DFF_X al_269819b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[10]));
  AL_DFF_X al_c748bb6f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[11]));
  AL_DFF_X al_6296777c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[12]));
  AL_DFF_X al_ae1847de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[13]));
  AL_DFF_X al_9626c91a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[14]));
  AL_DFF_X al_2d7b80c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[15]));
  AL_DFF_X al_390ef67f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[16]));
  AL_DFF_X al_c036586 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[17]));
  AL_DFF_X al_a78b54ea (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[18]));
  AL_DFF_X al_ec95e83d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[1]));
  AL_DFF_X al_c7621ed2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[19]));
  AL_DFF_X al_8d3f8651 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[20]));
  AL_DFF_X al_1475e152 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[21]));
  AL_DFF_X al_f798559e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[22]));
  AL_DFF_X al_bf1d07f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[23]));
  AL_DFF_X al_6e33e0e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[24]));
  AL_DFF_X al_15c0e11e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[25]));
  AL_DFF_X al_56a239db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[26]));
  AL_DFF_X al_930674c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[27]));
  AL_DFF_X al_d7e9be6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[28]));
  AL_DFF_X al_d59f556a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[2]));
  AL_DFF_X al_83f0e9b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[29]));
  AL_DFF_X al_bd5982ba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[30]));
  AL_DFF_X al_672f9309 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[31]));
  AL_DFF_X al_fc6e3acc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[32]));
  AL_DFF_X al_d8f77e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[33]));
  AL_DFF_X al_4feee2fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[34]));
  AL_DFF_X al_e4665d9f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[35]));
  AL_DFF_X al_16649cd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[36]));
  AL_DFF_X al_ffc2c867 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[37]));
  AL_DFF_X al_f015d31d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[38]));
  AL_DFF_X al_5c007dd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[3]));
  AL_DFF_X al_da9216c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[39]));
  AL_DFF_X al_66cf885e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[40]));
  AL_DFF_X al_18c8bac2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[41]));
  AL_DFF_X al_bccd2f0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[42]));
  AL_DFF_X al_c621c681 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[43]));
  AL_DFF_X al_44eb231a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[44]));
  AL_DFF_X al_1df9f81d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[45]));
  AL_DFF_X al_8f85a86d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[46]));
  AL_DFF_X al_bf3d95a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[47]));
  AL_DFF_X al_2ae9a81c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[4]));
  AL_DFF_X al_7f5213b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[5]));
  AL_DFF_X al_2b465c98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[6]));
  AL_DFF_X al_f02f6fe2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[7]));
  AL_DFF_X al_1ca6e0c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59124752[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3b63a678[8]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ea897437 (
    .a(al_8f041238[7]),
    .b(al_ac1cba4d[7]),
    .c(al_93915853),
    .o({al_6abbbc54,al_42247ac7[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_78561ff8 (
    .a(al_8f041238[8]),
    .b(al_ac1cba4d[8]),
    .c(al_6abbbc54),
    .o({al_aa70c10f,al_42247ac7[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fa02e757 (
    .a(al_8f041238[9]),
    .b(al_ac1cba4d[9]),
    .c(al_aa70c10f),
    .o({al_41b2a88c,al_42247ac7[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bfd8b692 (
    .a(al_8f041238[10]),
    .b(al_ac1cba4d[10]),
    .c(al_41b2a88c),
    .o({al_dde17c7f,al_42247ac7[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ef569ff3 (
    .a(al_8f041238[11]),
    .b(al_ac1cba4d[11]),
    .c(al_dde17c7f),
    .o({al_6df879f,al_42247ac7[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b91ad6b6 (
    .a(al_8f041238[12]),
    .b(al_ac1cba4d[12]),
    .c(al_6df879f),
    .o({al_ca3af73f,al_42247ac7[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4847f2f2 (
    .a(al_8f041238[13]),
    .b(al_ac1cba4d[13]),
    .c(al_ca3af73f),
    .o({al_b8b96eac,al_42247ac7[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f949f5f3 (
    .a(al_8f041238[14]),
    .b(al_ac1cba4d[14]),
    .c(al_b8b96eac),
    .o({al_d7300a25,al_42247ac7[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4607f45e (
    .a(al_8f041238[15]),
    .b(al_ac1cba4d[15]),
    .c(al_d7300a25),
    .o({al_9c595c5,al_42247ac7[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e4fd6652 (
    .a(al_8f041238[16]),
    .b(al_ac1cba4d[16]),
    .c(al_9c595c5),
    .o({al_b47bbe21,al_42247ac7[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_f4af5624 (
    .a(1'b0),
    .o({al_4e2c20db,open_n207}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_715bac1f (
    .a(al_8f041238[17]),
    .b(al_ac1cba4d[17]),
    .c(al_b47bbe21),
    .o({al_e295dc49,al_42247ac7[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f503564 (
    .a(al_8f041238[18]),
    .b(al_ac1cba4d[18]),
    .c(al_e295dc49),
    .o({al_85e166c5,al_42247ac7[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_963fc8b6 (
    .a(al_8f041238[19]),
    .b(al_ac1cba4d[19]),
    .c(al_85e166c5),
    .o({al_689afff7,al_42247ac7[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f9e50871 (
    .a(al_8f041238[20]),
    .b(al_ac1cba4d[20]),
    .c(al_689afff7),
    .o({al_36c0ab0e,al_42247ac7[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_41a7a67 (
    .a(al_8f041238[21]),
    .b(al_ac1cba4d[21]),
    .c(al_36c0ab0e),
    .o({al_9cf8f60d,al_42247ac7[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_374ee91d (
    .a(al_8f041238[22]),
    .b(al_ac1cba4d[22]),
    .c(al_9cf8f60d),
    .o({al_a8352957,al_42247ac7[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_68eab474 (
    .a(al_8f041238[23]),
    .b(al_ac1cba4d[23]),
    .c(al_a8352957),
    .o({al_be007839,al_42247ac7[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_870d76c3 (
    .a(al_8f041238[24]),
    .b(al_ac1cba4d[24]),
    .c(al_be007839),
    .o({al_66995ad4,al_42247ac7[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bc1ab4df (
    .a(al_8f041238[25]),
    .b(al_ac1cba4d[25]),
    .c(al_66995ad4),
    .o({al_4dcb599e,al_42247ac7[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5b4d67d9 (
    .a(al_8f041238[26]),
    .b(al_ac1cba4d[26]),
    .c(al_4dcb599e),
    .o({al_155419a5,al_42247ac7[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7a8aca0 (
    .a(al_8f041238[0]),
    .b(al_ac1cba4d[0]),
    .c(al_4e2c20db),
    .o({al_5334aacc,al_42247ac7[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_feee767e (
    .a(al_8f041238[27]),
    .b(al_ac1cba4d[27]),
    .c(al_155419a5),
    .o({al_49b8db26,al_42247ac7[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_5bcba84a (
    .a(al_8f041238[28]),
    .b(al_ac1cba4d[28]),
    .c(al_49b8db26),
    .o({al_8468641,al_42247ac7[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2938ffcf (
    .a(al_8f041238[29]),
    .b(al_ac1cba4d[29]),
    .c(al_8468641),
    .o({al_9f4fbb79,al_42247ac7[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4b0e5b1c (
    .a(al_8f041238[30]),
    .b(al_ac1cba4d[30]),
    .c(al_9f4fbb79),
    .o({al_732042af,al_42247ac7[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2fe82627 (
    .a(al_8f041238[31]),
    .b(al_ac1cba4d[31]),
    .c(al_732042af),
    .o({al_cd055708,al_42247ac7[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2f42e9fd (
    .a(al_8f041238[32]),
    .b(1'b0),
    .c(al_cd055708),
    .o({al_2e4b86ef,open_n208}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f5cbbe3f (
    .a(1'b0),
    .b(1'b1),
    .c(al_2e4b86ef),
    .o({open_n209,al_b84db2a6}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_efcb06dc (
    .a(al_8f041238[1]),
    .b(al_ac1cba4d[1]),
    .c(al_5334aacc),
    .o({al_c6f75c3f,al_42247ac7[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b7b591e8 (
    .a(al_8f041238[2]),
    .b(al_ac1cba4d[2]),
    .c(al_c6f75c3f),
    .o({al_d26c1ceb,al_42247ac7[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2c1cf3e0 (
    .a(al_8f041238[3]),
    .b(al_ac1cba4d[3]),
    .c(al_d26c1ceb),
    .o({al_22bff0ea,al_42247ac7[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f862e417 (
    .a(al_8f041238[4]),
    .b(al_ac1cba4d[4]),
    .c(al_22bff0ea),
    .o({al_38e51a5b,al_42247ac7[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2ea1b7d (
    .a(al_8f041238[5]),
    .b(al_ac1cba4d[5]),
    .c(al_38e51a5b),
    .o({al_6b77e7f1,al_42247ac7[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d6086ff2 (
    .a(al_8f041238[6]),
    .b(al_ac1cba4d[6]),
    .c(al_6b77e7f1),
    .o({al_93915853,al_42247ac7[6]}));
  AL_DFF_X al_c5b4f0ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f336c405[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f23786d8[0]));
  AL_DFF_X al_f24fa23e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[42]));
  AL_DFF_X al_b9510f91 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[43]));
  AL_DFF_X al_20066f77 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[44]));
  AL_DFF_X al_1ca1c8a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[45]));
  AL_DFF_X al_106f8dd8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[46]));
  AL_DFF_X al_a8b71ae8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[47]));
  AL_DFF_X al_cbc5759e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[48]));
  AL_DFF_X al_7cb801b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[49]));
  AL_DFF_X al_511f8172 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[50]));
  AL_DFF_X al_57e1bf3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[51]));
  AL_DFF_X al_a66c12b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[52]));
  AL_DFF_X al_31e45cb7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[53]));
  AL_DFF_X al_7c085f8e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[54]));
  AL_DFF_X al_92c4b746 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[55]));
  AL_DFF_X al_8c2dad86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[56]));
  AL_DFF_X al_a588634 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[57]));
  AL_DFF_X al_d5871ce6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[58]));
  AL_DFF_X al_d90784d7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[59]));
  AL_DFF_X al_bf6ed91a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[60]));
  AL_DFF_X al_56d1c28c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[61]));
  AL_DFF_X al_dc62cfbe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[62]));
  AL_DFF_X al_367e678b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[63]));
  AL_DFF_X al_6bd4ee74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[64]));
  AL_DFF_X al_6f2ed6f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[65]));
  AL_DFF_X al_57365eb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[66]));
  AL_DFF_X al_281ce4c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[67]));
  AL_DFF_X al_40217ef0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[68]));
  AL_DFF_X al_aeb72098 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[69]));
  AL_DFF_X al_ea50b466 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[70]));
  AL_DFF_X al_7e80172d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[71]));
  AL_DFF_X al_df8fdbed (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[72]));
  AL_DFF_X al_7b38333a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_28202fa7[74]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_68bb3ebd[73]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    al_de175db (
    .a(al_9459711),
    .b(al_57ac52e7),
    .o(al_41ebf214));
  AL_MAP_LUT6 #(
    .EQN("(~(B)*~(C)*~((~D*A))*~(E)*~(F)+~(B)*~(C)*~((~D*A))*E*~(F)+B*~(C)*~((~D*A))*E*~(F)+~(B)*~(C)*(~D*A)*E*~(F)+~(B)*~(C)*~((~D*A))*~(E)*F+B*~(C)*~((~D*A))*~(E)*F+~(B)*C*~((~D*A))*~(E)*F+~(B)*~(C)*(~D*A)*~(E)*F+B*~(C)*(~D*A)*~(E)*F+~(B)*~(C)*~((~D*A))*E*F+B*~(C)*~((~D*A))*E*F+~(B)*C*~((~D*A))*E*F+B*C*~((~D*A))*E*F+~(B)*~(C)*(~D*A)*E*F+B*~(C)*(~D*A)*E*F+~(B)*C*(~D*A)*E*F)"),
    .INIT(64'hff7f3f1f0f070301))
    al_d8b7d5de (
    .a(al_28202fa7[43]),
    .b(al_28202fa7[44]),
    .c(al_28202fa7[45]),
    .d(al_1d4399b1[43]),
    .e(al_1d4399b1[44]),
    .f(al_1d4399b1[45]),
    .o(al_526f98e2));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    al_6770bbdd (
    .a(al_1fb17bb2),
    .b(al_35fbae96),
    .c(al_453ca3a4),
    .o(al_e907e498));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_db31256b (
    .a(al_28202fa7[61]),
    .b(al_28202fa7[62]),
    .c(al_28202fa7[65]),
    .d(al_28202fa7[66]),
    .e(al_28202fa7[68]),
    .f(al_28202fa7[71]),
    .o(al_e1852c9f));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_2cf103f6 (
    .a(al_28202fa7[49]),
    .b(al_28202fa7[50]),
    .c(al_28202fa7[52]),
    .d(al_28202fa7[55]),
    .e(al_28202fa7[56]),
    .f(al_28202fa7[59]),
    .o(al_3432ca06));
  AL_MAP_LUT6 #(
    .EQN("(F@(E*D*C*B*~A))"),
    .INIT(64'hbfffffff40000000))
    al_9c07658d (
    .a(al_9459711),
    .b(al_e907e498),
    .c(al_e1852c9f),
    .d(al_3432ca06),
    .e(al_28202fa7[43]),
    .f(al_1d4399b1[43]),
    .o(al_7a8c14f1[43]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*C*D*E)"),
    .INIT(32'h40d0f4fd))
    al_6b8d7338 (
    .a(al_526f98e2),
    .b(al_28202fa7[46]),
    .c(al_28202fa7[47]),
    .d(al_1d4399b1[46]),
    .e(al_1d4399b1[47]),
    .o(al_9459711));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_6013e167 (
    .a(al_28202fa7[64]),
    .b(al_28202fa7[67]),
    .c(al_28202fa7[69]),
    .d(al_28202fa7[70]),
    .e(al_28202fa7[72]),
    .f(al_28202fa7[73]),
    .o(al_1fb17bb2));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_db5db90d (
    .a(al_28202fa7[53]),
    .b(al_28202fa7[54]),
    .c(al_28202fa7[57]),
    .d(al_28202fa7[58]),
    .e(al_28202fa7[60]),
    .f(al_28202fa7[63]),
    .o(al_35fbae96));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_9689c7d7 (
    .a(al_28202fa7[48]),
    .b(al_28202fa7[51]),
    .c(al_28202fa7[74]),
    .o(al_453ca3a4));
  AL_MAP_LUT5 #(
    .EQN("(B*A*(D@(~E*C)))"),
    .INIT(32'h88000880))
    al_62a0a41d (
    .a(al_e1852c9f),
    .b(al_3432ca06),
    .c(al_28202fa7[43]),
    .d(al_28202fa7[44]),
    .e(al_1d4399b1[43]),
    .o(al_5b27964b));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*B*~A))"),
    .INIT(16'hbf40))
    al_cf17b53d (
    .a(al_9459711),
    .b(al_e907e498),
    .c(al_5b27964b),
    .d(al_1d4399b1[44]),
    .o(al_7a8c14f1[44]));
  AL_MAP_LUT5 #(
    .EQN("(C@(B*~((~D*A))*~(E)+~(B)*(~D*A)*~(E)+B*(~D*A)*~(E)+B*(~D*A)*E))"),
    .INIT(32'hf0783c1e))
    al_715d55f4 (
    .a(al_28202fa7[43]),
    .b(al_28202fa7[44]),
    .c(al_28202fa7[45]),
    .d(al_1d4399b1[43]),
    .e(al_1d4399b1[44]),
    .o(al_e6e3fffa));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*B*~A))"),
    .INIT(16'hbf40))
    al_7076dd84 (
    .a(al_9459711),
    .b(al_57ac52e7),
    .c(al_e6e3fffa),
    .d(al_1d4399b1[45]),
    .o(al_7a8c14f1[45]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_6340aaa7 (
    .a(al_1fb17bb2),
    .b(al_35fbae96),
    .c(al_453ca3a4),
    .d(al_e1852c9f),
    .e(al_3432ca06),
    .o(al_57ac52e7));
  AL_MAP_LUT5 #(
    .EQN("(E@(B*~A*~(D@C)))"),
    .INIT(32'hbffb4004))
    al_ce04fd1e (
    .a(al_9459711),
    .b(al_57ac52e7),
    .c(al_526f98e2),
    .d(al_28202fa7[46]),
    .e(al_1d4399b1[46]),
    .o(al_7a8c14f1[46]));
  AL_MAP_LUT6 #(
    .EQN("(F*~(A*~(D@(B*~(C)*~(E)+~(B)*~(C)*E+B*~(C)*E+B*C*E))))"),
    .INIT(64'h75dff75d00000000))
    al_c42bbb1 (
    .a(al_57ac52e7),
    .b(al_526f98e2),
    .c(al_28202fa7[46]),
    .d(al_28202fa7[47]),
    .e(al_1d4399b1[46]),
    .f(al_1d4399b1[47]),
    .o(al_7a8c14f1[47]));
  AL_DFF_X al_67624b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[0]));
  AL_DFF_X al_c3a708d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[9]));
  AL_DFF_X al_43ffedde (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[10]));
  AL_DFF_X al_9e6730d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[11]));
  AL_DFF_X al_d1b3e088 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[12]));
  AL_DFF_X al_ffbede16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[13]));
  AL_DFF_X al_aa788c7f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[14]));
  AL_DFF_X al_4728c2a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[15]));
  AL_DFF_X al_2cd37b08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[16]));
  AL_DFF_X al_216e4c19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[17]));
  AL_DFF_X al_16b6cedb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[18]));
  AL_DFF_X al_9386a037 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[1]));
  AL_DFF_X al_4859d7c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[19]));
  AL_DFF_X al_dfd0e35b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[20]));
  AL_DFF_X al_13e99445 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[21]));
  AL_DFF_X al_3d8d32b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[22]));
  AL_DFF_X al_148fbc01 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[23]));
  AL_DFF_X al_80ae70ab (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[24]));
  AL_DFF_X al_830ce8ce (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[25]));
  AL_DFF_X al_4f313285 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[26]));
  AL_DFF_X al_45947bf4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[27]));
  AL_DFF_X al_7571b095 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[28]));
  AL_DFF_X al_ab027576 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[2]));
  AL_DFF_X al_3c401e4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[29]));
  AL_DFF_X al_167df66a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[30]));
  AL_DFF_X al_b42f11ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[31]));
  AL_DFF_X al_14c37c8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[32]));
  AL_DFF_X al_5229687 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[33]));
  AL_DFF_X al_a61301c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[34]));
  AL_DFF_X al_7e65217d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[35]));
  AL_DFF_X al_395f7bdc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[36]));
  AL_DFF_X al_70f8d71 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[37]));
  AL_DFF_X al_b44a1705 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[38]));
  AL_DFF_X al_adbe07f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[3]));
  AL_DFF_X al_8080d80f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[39]));
  AL_DFF_X al_a69bf41d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[40]));
  AL_DFF_X al_7e2f9709 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[41]));
  AL_DFF_X al_542c3a1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[42]));
  AL_DFF_X al_a452b498 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[43]));
  AL_DFF_X al_1995e75e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[44]));
  AL_DFF_X al_916ce359 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[45]));
  AL_DFF_X al_49f68f85 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[46]));
  AL_DFF_X al_9b506140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7a8c14f1[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[47]));
  AL_DFF_X al_fb760e2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[4]));
  AL_DFF_X al_2700ec19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[5]));
  AL_DFF_X al_fdbdef28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[6]));
  AL_DFF_X al_8fbbae9d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[7]));
  AL_DFF_X al_4423c666 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1d4399b1[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_1b3e91c5[8]));
  AL_DFF_X al_60368985 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_41ebf214),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[0]));
  AL_DFF_X al_c5f86dd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_917df14b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[1]));
  AL_DFF_X al_9ccf400 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_917df14b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[2]));
  AL_DFF_X al_d7435a14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_917df14b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[3]));
  AL_DFF_X al_5321d04b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_917df14b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4682e2e2[4]));
  AL_DFF_X al_d0c29a4f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f23786d8[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6e4d5f5f[0]));
  AL_DFF_X al_bbdbda09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[41]));
  AL_DFF_X al_b4017ff (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[42]));
  AL_DFF_X al_ab4f4118 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[43]));
  AL_DFF_X al_296f6990 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[44]));
  AL_DFF_X al_671979a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[45]));
  AL_DFF_X al_acd2e2fd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[46]));
  AL_DFF_X al_581df90b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[47]));
  AL_DFF_X al_1abe2e36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[48]));
  AL_DFF_X al_154bfdd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[49]));
  AL_DFF_X al_46b10b4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[50]));
  AL_DFF_X al_aa0e753 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[51]));
  AL_DFF_X al_83ecf292 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[52]));
  AL_DFF_X al_fa34fcc8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[53]));
  AL_DFF_X al_5001d0c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[54]));
  AL_DFF_X al_2ba5074a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[55]));
  AL_DFF_X al_a3e25a44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[56]));
  AL_DFF_X al_a5b864fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[57]));
  AL_DFF_X al_11f6def3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[58]));
  AL_DFF_X al_3614f507 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[59]));
  AL_DFF_X al_6b62cc8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[60]));
  AL_DFF_X al_95684a09 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[61]));
  AL_DFF_X al_207c3aad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[62]));
  AL_DFF_X al_7b133c8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[63]));
  AL_DFF_X al_1f7dba22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[64]));
  AL_DFF_X al_ac9b783d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[65]));
  AL_DFF_X al_3681bea2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[66]));
  AL_DFF_X al_d714f156 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[67]));
  AL_DFF_X al_512cc40e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[68]));
  AL_DFF_X al_60b081a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[69]));
  AL_DFF_X al_708b29e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[70]));
  AL_DFF_X al_9cd7c324 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[71]));
  AL_DFF_X al_d832a4a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_68bb3ebd[73]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2a9de02[72]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_bc993dfd (
    .a(1'b0),
    .o({al_2b438376,open_n212}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_b57ea34e (
    .a(al_1b3e91c5[42]),
    .b(al_68bb3ebd[42]),
    .c(al_2b438376),
    .o({al_ca3e9bc8,al_504aeee4[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_767558c6 (
    .a(al_1b3e91c5[43]),
    .b(al_68bb3ebd[43]),
    .c(al_ca3e9bc8),
    .o({al_464b5ec,al_504aeee4[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7b9955b (
    .a(al_1b3e91c5[44]),
    .b(al_68bb3ebd[44]),
    .c(al_464b5ec),
    .o({al_a0e81a0c,al_504aeee4[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9bd0f4ac (
    .a(al_1b3e91c5[45]),
    .b(al_68bb3ebd[45]),
    .c(al_a0e81a0c),
    .o({al_6e619896,al_504aeee4[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_76c7052b (
    .a(al_1b3e91c5[46]),
    .b(al_68bb3ebd[46]),
    .c(al_6e619896),
    .o({al_f3664844,al_504aeee4[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d497567a (
    .a(al_1b3e91c5[47]),
    .b(al_68bb3ebd[47]),
    .c(al_f3664844),
    .o({al_eb180f53,al_504aeee4[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_17cb9dc2 (
    .c(al_eb180f53),
    .o({open_n215,al_504aeee4[6]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d5573861 (
    .a(al_b9439b67),
    .b(al_1b3e91c5[42]),
    .c(al_504aeee4[0]),
    .o(al_7d7cdb8e[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cd3e798f (
    .a(al_b9439b67),
    .b(al_1b3e91c5[43]),
    .c(al_504aeee4[1]),
    .o(al_7d7cdb8e[43]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_7dd115d (
    .a(al_68bb3ebd[68]),
    .b(al_68bb3ebd[69]),
    .c(al_68bb3ebd[70]),
    .d(al_68bb3ebd[71]),
    .e(al_68bb3ebd[72]),
    .f(al_68bb3ebd[73]),
    .o(al_ad51aadd));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    al_4a753f19 (
    .a(al_ad51aadd),
    .b(al_aa6720b4),
    .c(al_82c92bf1),
    .d(al_51ccac31),
    .e(al_a50d3ef5),
    .o(al_b9439b67));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6d7321a7 (
    .a(al_b9439b67),
    .b(al_1b3e91c5[44]),
    .c(al_504aeee4[2]),
    .o(al_7d7cdb8e[44]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_772a56ff (
    .a(al_68bb3ebd[62]),
    .b(al_68bb3ebd[63]),
    .c(al_68bb3ebd[64]),
    .d(al_68bb3ebd[65]),
    .e(al_68bb3ebd[66]),
    .f(al_68bb3ebd[67]),
    .o(al_aa6720b4));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_9cb786f7 (
    .a(al_68bb3ebd[56]),
    .b(al_68bb3ebd[57]),
    .c(al_68bb3ebd[58]),
    .d(al_68bb3ebd[59]),
    .e(al_68bb3ebd[60]),
    .f(al_68bb3ebd[61]),
    .o(al_82c92bf1));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_f3036be8 (
    .a(al_68bb3ebd[50]),
    .b(al_68bb3ebd[51]),
    .c(al_68bb3ebd[52]),
    .d(al_68bb3ebd[53]),
    .e(al_68bb3ebd[54]),
    .f(al_68bb3ebd[55]),
    .o(al_51ccac31));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    al_bb2cc98 (
    .a(al_68bb3ebd[48]),
    .b(al_68bb3ebd[49]),
    .c(al_504aeee4[6]),
    .o(al_a50d3ef5));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f380b667 (
    .a(al_b9439b67),
    .b(al_1b3e91c5[45]),
    .c(al_504aeee4[3]),
    .o(al_7d7cdb8e[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_8ac7c6d0 (
    .a(al_b9439b67),
    .b(al_1b3e91c5[46]),
    .c(al_504aeee4[4]),
    .o(al_7d7cdb8e[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6a6ea6ae (
    .a(al_b9439b67),
    .b(al_1b3e91c5[47]),
    .c(al_504aeee4[5]),
    .o(al_7d7cdb8e[47]));
  AL_DFF_X al_69dfe244 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[0]));
  AL_DFF_X al_aa24be8d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[9]));
  AL_DFF_X al_34670a3b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[10]));
  AL_DFF_X al_9cec3d2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[11]));
  AL_DFF_X al_8f6b2215 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[12]));
  AL_DFF_X al_e84c9f27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[13]));
  AL_DFF_X al_5e110ec2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[14]));
  AL_DFF_X al_4f51cabe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[15]));
  AL_DFF_X al_4e65cdc9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[16]));
  AL_DFF_X al_44f1e012 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[17]));
  AL_DFF_X al_29f2edee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[18]));
  AL_DFF_X al_885213f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[1]));
  AL_DFF_X al_7c65b883 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[19]));
  AL_DFF_X al_4c5f209b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[20]));
  AL_DFF_X al_2c4f00f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[21]));
  AL_DFF_X al_c5f4e4b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[22]));
  AL_DFF_X al_b256e95c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[23]));
  AL_DFF_X al_86397550 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[24]));
  AL_DFF_X al_d8d511a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[25]));
  AL_DFF_X al_2c02df3e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[26]));
  AL_DFF_X al_b258723a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[27]));
  AL_DFF_X al_bbf1c243 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[28]));
  AL_DFF_X al_6f37bca4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[2]));
  AL_DFF_X al_97ded0fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[29]));
  AL_DFF_X al_f85b5c89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[30]));
  AL_DFF_X al_e3a3581b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[31]));
  AL_DFF_X al_1ff1bc82 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[32]));
  AL_DFF_X al_82a490dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[33]));
  AL_DFF_X al_8dadb241 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[34]));
  AL_DFF_X al_5c2db451 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[35]));
  AL_DFF_X al_892af1e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[36]));
  AL_DFF_X al_bf8d575b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[37]));
  AL_DFF_X al_86855c36 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[38]));
  AL_DFF_X al_fec29d24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[3]));
  AL_DFF_X al_a2a4422b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[39]));
  AL_DFF_X al_8f1643d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[40]));
  AL_DFF_X al_95b91672 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[41]));
  AL_DFF_X al_4eb3167e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[42]));
  AL_DFF_X al_936d0732 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[43]));
  AL_DFF_X al_62c21e25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[44]));
  AL_DFF_X al_4f5923c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[45]));
  AL_DFF_X al_b56684db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[46]));
  AL_DFF_X al_c93ca04d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_7d7cdb8e[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[47]));
  AL_DFF_X al_136526d0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[4]));
  AL_DFF_X al_5dc72afd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[5]));
  AL_DFF_X al_f54fda76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[6]));
  AL_DFF_X al_b5c387a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[7]));
  AL_DFF_X al_1f16b017 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1b3e91c5[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_15503509[8]));
  AL_DFF_X al_6d4e73a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_b9439b67),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[0]));
  AL_DFF_X al_737090bb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[1]));
  AL_DFF_X al_45abfbf5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[2]));
  AL_DFF_X al_18e7b7a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[3]));
  AL_DFF_X al_bb26e1fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[4]));
  AL_DFF_X al_8c7a490d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4682e2e2[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_22a22ff3[5]));
  AL_DFF_X al_f7f0d87b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_6e4d5f5f[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d255f877[0]));
  AL_DFF_X al_e77d71a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[40]));
  AL_DFF_X al_446faf0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[41]));
  AL_DFF_X al_3a3671e7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[42]));
  AL_DFF_X al_5102644d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[43]));
  AL_DFF_X al_c424a8d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[44]));
  AL_DFF_X al_e8da13e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[45]));
  AL_DFF_X al_ff2d169f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[46]));
  AL_DFF_X al_8fde187b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[47]));
  AL_DFF_X al_7419ade4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[48]));
  AL_DFF_X al_fe561575 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[49]));
  AL_DFF_X al_208aac98 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[50]));
  AL_DFF_X al_768521c5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[51]));
  AL_DFF_X al_29a54be7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[52]));
  AL_DFF_X al_973be54b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[53]));
  AL_DFF_X al_bbfe44a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[54]));
  AL_DFF_X al_f96eba52 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[55]));
  AL_DFF_X al_fba66cd1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[56]));
  AL_DFF_X al_fd2d0c1d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[57]));
  AL_DFF_X al_4992630 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[58]));
  AL_DFF_X al_ed8c9ce8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[59]));
  AL_DFF_X al_f51081a6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[60]));
  AL_DFF_X al_5d748987 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[61]));
  AL_DFF_X al_7a31da03 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[62]));
  AL_DFF_X al_d36dd1ee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[63]));
  AL_DFF_X al_cbc2439a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[64]));
  AL_DFF_X al_cdd1574c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[65]));
  AL_DFF_X al_f30db30d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[66]));
  AL_DFF_X al_ebdd36b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[67]));
  AL_DFF_X al_99328fad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[68]));
  AL_DFF_X al_275bd682 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[69]));
  AL_DFF_X al_ac26254b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[70]));
  AL_DFF_X al_1190754d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f2a9de02[72]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5206392b[71]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_ea7d4896 (
    .a(1'b0),
    .o({al_24f0c9b4,open_n218}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_15aa0ba7 (
    .a(al_15503509[41]),
    .b(al_f2a9de02[41]),
    .c(al_24f0c9b4),
    .o({al_8e479b1b,al_b9ac5fd4[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7c29e9dc (
    .a(al_15503509[42]),
    .b(al_f2a9de02[42]),
    .c(al_8e479b1b),
    .o({al_6aa12cb6,al_b9ac5fd4[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_180912c3 (
    .a(al_15503509[43]),
    .b(al_f2a9de02[43]),
    .c(al_6aa12cb6),
    .o({al_1d3f4f78,al_b9ac5fd4[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ddf981e2 (
    .a(al_15503509[44]),
    .b(al_f2a9de02[44]),
    .c(al_1d3f4f78),
    .o({al_63e4776,al_b9ac5fd4[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_beaef896 (
    .a(al_15503509[45]),
    .b(al_f2a9de02[45]),
    .c(al_63e4776),
    .o({al_fb5dab05,al_b9ac5fd4[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ff3f86f7 (
    .a(al_15503509[46]),
    .b(al_f2a9de02[46]),
    .c(al_fb5dab05),
    .o({al_2e3e139,al_b9ac5fd4[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3a6a9953 (
    .a(al_15503509[47]),
    .b(al_f2a9de02[47]),
    .c(al_2e3e139),
    .o({al_92d8d26e,al_b9ac5fd4[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_73d217cc (
    .c(al_92d8d26e),
    .o({open_n221,al_b9ac5fd4[7]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_c1d4c70e (
    .a(al_f2a9de02[68]),
    .b(al_f2a9de02[69]),
    .c(al_f2a9de02[70]),
    .d(al_f2a9de02[71]),
    .e(al_f2a9de02[72]),
    .f(al_b9ac5fd4[7]),
    .o(al_94cd12cf));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_32b70cba (
    .a(al_c1da9790),
    .b(al_15503509[41]),
    .c(al_b9ac5fd4[0]),
    .o(al_78306f09[41]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_d244d681 (
    .a(al_f2a9de02[62]),
    .b(al_f2a9de02[63]),
    .c(al_f2a9de02[64]),
    .d(al_f2a9de02[65]),
    .e(al_f2a9de02[66]),
    .f(al_f2a9de02[67]),
    .o(al_31ed294d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_5368fd1e (
    .a(al_f2a9de02[56]),
    .b(al_f2a9de02[57]),
    .c(al_f2a9de02[58]),
    .d(al_f2a9de02[59]),
    .e(al_f2a9de02[60]),
    .f(al_f2a9de02[61]),
    .o(al_58d02051));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_51cdcbf (
    .a(al_f2a9de02[50]),
    .b(al_f2a9de02[51]),
    .c(al_f2a9de02[52]),
    .d(al_f2a9de02[53]),
    .e(al_f2a9de02[54]),
    .f(al_f2a9de02[55]),
    .o(al_1024d4fd));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*D*C*B*A)"),
    .INIT(64'h0000000000008000))
    al_cd06b53b (
    .a(al_94cd12cf),
    .b(al_31ed294d),
    .c(al_58d02051),
    .d(al_1024d4fd),
    .e(al_f2a9de02[48]),
    .f(al_f2a9de02[49]),
    .o(al_c1da9790));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_47cd0b20 (
    .a(al_c1da9790),
    .b(al_15503509[42]),
    .c(al_b9ac5fd4[1]),
    .o(al_78306f09[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3f0380ee (
    .a(al_c1da9790),
    .b(al_15503509[43]),
    .c(al_b9ac5fd4[2]),
    .o(al_78306f09[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7dfb6c89 (
    .a(al_c1da9790),
    .b(al_15503509[44]),
    .c(al_b9ac5fd4[3]),
    .o(al_78306f09[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1ee8ea3a (
    .a(al_c1da9790),
    .b(al_15503509[45]),
    .c(al_b9ac5fd4[4]),
    .o(al_78306f09[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_f888c136 (
    .a(al_c1da9790),
    .b(al_15503509[46]),
    .c(al_b9ac5fd4[5]),
    .o(al_78306f09[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_a0e8cee7 (
    .a(al_c1da9790),
    .b(al_15503509[47]),
    .c(al_b9ac5fd4[6]),
    .o(al_78306f09[47]));
  AL_DFF_X al_4ff7d84a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[0]));
  AL_DFF_X al_cfdc3e17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[9]));
  AL_DFF_X al_97de1911 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[10]));
  AL_DFF_X al_7f02a4af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[11]));
  AL_DFF_X al_35a7a994 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[12]));
  AL_DFF_X al_38e84c27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[13]));
  AL_DFF_X al_e3be7404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[14]));
  AL_DFF_X al_44334c31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[15]));
  AL_DFF_X al_afa18a08 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[16]));
  AL_DFF_X al_78accdd2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[17]));
  AL_DFF_X al_909f496d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[18]));
  AL_DFF_X al_e64226eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[1]));
  AL_DFF_X al_b1298452 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[19]));
  AL_DFF_X al_6aef2061 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[20]));
  AL_DFF_X al_d2c5f6b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[21]));
  AL_DFF_X al_dc11ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[22]));
  AL_DFF_X al_2713b67e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[23]));
  AL_DFF_X al_62015d59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[24]));
  AL_DFF_X al_8fa4e871 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[25]));
  AL_DFF_X al_dfa8c073 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[26]));
  AL_DFF_X al_358dc259 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[27]));
  AL_DFF_X al_332bc2bf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[28]));
  AL_DFF_X al_780ccc0c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[2]));
  AL_DFF_X al_201ce062 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[29]));
  AL_DFF_X al_6f723813 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[30]));
  AL_DFF_X al_a4337ba0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[31]));
  AL_DFF_X al_c1d9154a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[32]));
  AL_DFF_X al_4ecae0c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[33]));
  AL_DFF_X al_d4763e5d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[34]));
  AL_DFF_X al_174d20cb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[35]));
  AL_DFF_X al_7cb06c9c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[36]));
  AL_DFF_X al_d2f22fee (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[37]));
  AL_DFF_X al_a373ee41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[38]));
  AL_DFF_X al_f241805c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[3]));
  AL_DFF_X al_4daae9af (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[39]));
  AL_DFF_X al_1d4d612d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[40]));
  AL_DFF_X al_7830bea8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[41]));
  AL_DFF_X al_37855439 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[42]));
  AL_DFF_X al_f7e07093 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[43]));
  AL_DFF_X al_de900bf9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[44]));
  AL_DFF_X al_d74f4d80 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[45]));
  AL_DFF_X al_cdef273 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[46]));
  AL_DFF_X al_9ff5483 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_78306f09[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[47]));
  AL_DFF_X al_ecfeb63a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[4]));
  AL_DFF_X al_911d6634 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[5]));
  AL_DFF_X al_8fdb9581 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[6]));
  AL_DFF_X al_9290b1df (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[7]));
  AL_DFF_X al_d9f92c15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_15503509[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_59bef53b[8]));
  AL_DFF_X al_61dc39c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1da9790),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[0]));
  AL_DFF_X al_b3f92f30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[1]));
  AL_DFF_X al_f1809f8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[2]));
  AL_DFF_X al_416f7ccf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[3]));
  AL_DFF_X al_f73f6fa5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[4]));
  AL_DFF_X al_7628f970 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[5]));
  AL_DFF_X al_4ee3f5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_22a22ff3[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9c3e2402[6]));
  AL_DFF_X al_c82698cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d255f877[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_30922aac[0]));
  AL_DFF_X al_ba344f29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[39]));
  AL_DFF_X al_5e85ba55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[40]));
  AL_DFF_X al_6ea0f290 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[41]));
  AL_DFF_X al_5bc50a00 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[42]));
  AL_DFF_X al_c1dbfdfc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[43]));
  AL_DFF_X al_18a1b86 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[44]));
  AL_DFF_X al_4cfe9dd9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[45]));
  AL_DFF_X al_71f5132d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[46]));
  AL_DFF_X al_e8d76e68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[47]));
  AL_DFF_X al_c0bdccae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[48]));
  AL_DFF_X al_6dff7a25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[49]));
  AL_DFF_X al_4abb60fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[50]));
  AL_DFF_X al_338673c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[51]));
  AL_DFF_X al_2b924789 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[52]));
  AL_DFF_X al_69271171 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[53]));
  AL_DFF_X al_f7f5c4b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[54]));
  AL_DFF_X al_3d717a6e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[55]));
  AL_DFF_X al_bcb69af1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[56]));
  AL_DFF_X al_c1367c2b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[57]));
  AL_DFF_X al_154c1d9a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[58]));
  AL_DFF_X al_159ed4cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[59]));
  AL_DFF_X al_b8c0c207 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[60]));
  AL_DFF_X al_9f321509 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[61]));
  AL_DFF_X al_b7035865 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[62]));
  AL_DFF_X al_934249b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[63]));
  AL_DFF_X al_f0aa6d4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[64]));
  AL_DFF_X al_c01904dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[65]));
  AL_DFF_X al_7c33b573 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[66]));
  AL_DFF_X al_b979a4e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[67]));
  AL_DFF_X al_bb21c38b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[68]));
  AL_DFF_X al_8ff98fc4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[69]));
  AL_DFF_X al_9225514d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5206392b[71]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_d6cb04b6[70]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_86bfeb89 (
    .a(1'b0),
    .o({al_6cad4dc9,open_n224}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_242792f6 (
    .a(al_59bef53b[40]),
    .b(al_5206392b[40]),
    .c(al_6cad4dc9),
    .o({al_2abe7dd5,al_f87eab88[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d8dd5e9f (
    .a(al_59bef53b[41]),
    .b(al_5206392b[41]),
    .c(al_2abe7dd5),
    .o({al_441d631,al_f87eab88[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_a07563d5 (
    .a(al_59bef53b[42]),
    .b(al_5206392b[42]),
    .c(al_441d631),
    .o({al_f3239c7d,al_f87eab88[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4c8a5b0b (
    .a(al_59bef53b[43]),
    .b(al_5206392b[43]),
    .c(al_f3239c7d),
    .o({al_b87907a9,al_f87eab88[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_60de78b1 (
    .a(al_59bef53b[44]),
    .b(al_5206392b[44]),
    .c(al_b87907a9),
    .o({al_90f0f7d8,al_f87eab88[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_8cbeafce (
    .a(al_59bef53b[45]),
    .b(al_5206392b[45]),
    .c(al_90f0f7d8),
    .o({al_a4b7f674,al_f87eab88[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_c1ca04a9 (
    .a(al_59bef53b[46]),
    .b(al_5206392b[46]),
    .c(al_a4b7f674),
    .o({al_7076449e,al_f87eab88[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_e4bef42b (
    .a(al_59bef53b[47]),
    .b(al_5206392b[47]),
    .c(al_7076449e),
    .o({al_8e44a4d6,al_f87eab88[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4774f25e (
    .c(al_8e44a4d6),
    .o({open_n227,al_f87eab88[8]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_560f3511 (
    .a(al_1881b524),
    .b(al_59bef53b[40]),
    .c(al_f87eab88[0]),
    .o(al_601b9c02[40]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_c86c70b6 (
    .a(al_5206392b[66]),
    .b(al_5206392b[67]),
    .c(al_5206392b[68]),
    .d(al_5206392b[69]),
    .e(al_5206392b[70]),
    .f(al_5206392b[71]),
    .o(al_4ff3fb03));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_2751844f (
    .a(al_1881b524),
    .b(al_59bef53b[41]),
    .c(al_f87eab88[1]),
    .o(al_601b9c02[41]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_4971210f (
    .a(al_5206392b[60]),
    .b(al_5206392b[61]),
    .c(al_5206392b[62]),
    .d(al_5206392b[63]),
    .e(al_5206392b[64]),
    .f(al_5206392b[65]),
    .o(al_724c9346));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_c63fb61c (
    .a(al_5206392b[54]),
    .b(al_5206392b[55]),
    .c(al_5206392b[56]),
    .d(al_5206392b[57]),
    .e(al_5206392b[58]),
    .f(al_5206392b[59]),
    .o(al_654ec6c7));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_161c873e (
    .a(al_5206392b[48]),
    .b(al_5206392b[49]),
    .c(al_5206392b[50]),
    .d(al_5206392b[51]),
    .e(al_5206392b[52]),
    .f(al_5206392b[53]),
    .o(al_db43acf6));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    al_d678e241 (
    .a(al_4ff3fb03),
    .b(al_724c9346),
    .c(al_654ec6c7),
    .d(al_db43acf6),
    .e(al_f87eab88[8]),
    .o(al_1881b524));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ad4d8f76 (
    .a(al_1881b524),
    .b(al_59bef53b[42]),
    .c(al_f87eab88[2]),
    .o(al_601b9c02[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_16af9e6f (
    .a(al_1881b524),
    .b(al_59bef53b[43]),
    .c(al_f87eab88[3]),
    .o(al_601b9c02[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1308b02c (
    .a(al_1881b524),
    .b(al_59bef53b[44]),
    .c(al_f87eab88[4]),
    .o(al_601b9c02[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_94c8cdc7 (
    .a(al_1881b524),
    .b(al_59bef53b[45]),
    .c(al_f87eab88[5]),
    .o(al_601b9c02[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_9cc9c7bc (
    .a(al_1881b524),
    .b(al_59bef53b[46]),
    .c(al_f87eab88[6]),
    .o(al_601b9c02[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ea4fe816 (
    .a(al_1881b524),
    .b(al_59bef53b[47]),
    .c(al_f87eab88[7]),
    .o(al_601b9c02[47]));
  AL_DFF_X al_fb22c32 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[0]));
  AL_DFF_X al_8c6b9882 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[9]));
  AL_DFF_X al_706b48d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[10]));
  AL_DFF_X al_bcd366fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[11]));
  AL_DFF_X al_af535c2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[12]));
  AL_DFF_X al_f7377aa1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[13]));
  AL_DFF_X al_92b03dca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[14]));
  AL_DFF_X al_23c6e620 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[15]));
  AL_DFF_X al_4627cc84 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[16]));
  AL_DFF_X al_9f364fe7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[17]));
  AL_DFF_X al_76eece0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[18]));
  AL_DFF_X al_ab07a2a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[1]));
  AL_DFF_X al_7cbc43c9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[19]));
  AL_DFF_X al_1502f910 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[20]));
  AL_DFF_X al_22b95b40 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[21]));
  AL_DFF_X al_34ee9d2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[22]));
  AL_DFF_X al_c529f40a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[23]));
  AL_DFF_X al_f90e4146 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[24]));
  AL_DFF_X al_266160fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[25]));
  AL_DFF_X al_f9488d30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[26]));
  AL_DFF_X al_506f2cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[27]));
  AL_DFF_X al_d5b0ce59 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[28]));
  AL_DFF_X al_ffe0e404 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[2]));
  AL_DFF_X al_3f6c1bd0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[29]));
  AL_DFF_X al_7743774a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[30]));
  AL_DFF_X al_2367aa20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[31]));
  AL_DFF_X al_6ef77cc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[32]));
  AL_DFF_X al_9b369669 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[33]));
  AL_DFF_X al_75055aba (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[34]));
  AL_DFF_X al_5c9a90e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[35]));
  AL_DFF_X al_89a75d6a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[36]));
  AL_DFF_X al_ef99cf3a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[37]));
  AL_DFF_X al_245dae74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[38]));
  AL_DFF_X al_21cf5cc0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[3]));
  AL_DFF_X al_89347f42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[39]));
  AL_DFF_X al_1209e91f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[40]));
  AL_DFF_X al_db3f12e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[41]));
  AL_DFF_X al_30d27b44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[42]));
  AL_DFF_X al_15f2f1c6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[43]));
  AL_DFF_X al_754c0140 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[44]));
  AL_DFF_X al_63901767 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[45]));
  AL_DFF_X al_c7fe6c5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[46]));
  AL_DFF_X al_50e5e56c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_601b9c02[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[47]));
  AL_DFF_X al_d5c56dbf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[4]));
  AL_DFF_X al_5aae32d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[5]));
  AL_DFF_X al_5177f848 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[6]));
  AL_DFF_X al_8e34ae55 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[7]));
  AL_DFF_X al_1665c65d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_59bef53b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f7a9a92b[8]));
  AL_DFF_X al_9bb3eb50 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_1881b524),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[0]));
  AL_DFF_X al_c5cd1544 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[1]));
  AL_DFF_X al_c84db15d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[2]));
  AL_DFF_X al_7b220268 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[3]));
  AL_DFF_X al_709e9629 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[4]));
  AL_DFF_X al_65175b92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[5]));
  AL_DFF_X al_5591c387 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[6]));
  AL_DFF_X al_ed963c22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_9c3e2402[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4dd3fb65[7]));
  AL_DFF_X al_fb7eed2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_30922aac[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_36d845bb[0]));
  AL_DFF_X al_546a979f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[38]));
  AL_DFF_X al_4af8b9a4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[39]));
  AL_DFF_X al_797a2d65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[40]));
  AL_DFF_X al_d608e00d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[41]));
  AL_DFF_X al_d90dba44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[42]));
  AL_DFF_X al_89e9f626 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[43]));
  AL_DFF_X al_129ca994 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[44]));
  AL_DFF_X al_f48eabd4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[45]));
  AL_DFF_X al_e3b61b4e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[46]));
  AL_DFF_X al_af7b09de (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[47]));
  AL_DFF_X al_25a5df5a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[48]));
  AL_DFF_X al_90af9f48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[49]));
  AL_DFF_X al_9b97099e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[50]));
  AL_DFF_X al_a178b03a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[51]));
  AL_DFF_X al_fedd492b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[52]));
  AL_DFF_X al_ca5f9de5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[53]));
  AL_DFF_X al_b5096629 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[54]));
  AL_DFF_X al_3549bac8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[55]));
  AL_DFF_X al_edeabf2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[56]));
  AL_DFF_X al_90e09490 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[57]));
  AL_DFF_X al_4fd0e29d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[58]));
  AL_DFF_X al_7dd6e2e1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[59]));
  AL_DFF_X al_8b6476d9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[60]));
  AL_DFF_X al_eb5ae236 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[61]));
  AL_DFF_X al_af9a20b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[62]));
  AL_DFF_X al_bc13fa94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[63]));
  AL_DFF_X al_fe7624cd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[64]));
  AL_DFF_X al_225430fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[65]));
  AL_DFF_X al_aaa60b94 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[66]));
  AL_DFF_X al_8e91b8fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[67]));
  AL_DFF_X al_75108b05 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[68]));
  AL_DFF_X al_c59aed8c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_d6cb04b6[70]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_c1960abd[69]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_5adae02f (
    .a(1'b0),
    .o({al_ee4e9a87,open_n230}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_23275c4a (
    .a(al_f7a9a92b[39]),
    .b(al_d6cb04b6[39]),
    .c(al_ee4e9a87),
    .o({al_ea6aa5ed,al_5b8748c3[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_3c89d57c (
    .a(al_f7a9a92b[40]),
    .b(al_d6cb04b6[40]),
    .c(al_ea6aa5ed),
    .o({al_d4f16200,al_5b8748c3[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_af058505 (
    .a(al_f7a9a92b[41]),
    .b(al_d6cb04b6[41]),
    .c(al_d4f16200),
    .o({al_ee99ca7f,al_5b8748c3[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_1c856914 (
    .a(al_f7a9a92b[42]),
    .b(al_d6cb04b6[42]),
    .c(al_ee99ca7f),
    .o({al_b8f391da,al_5b8748c3[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fc2c9df9 (
    .a(al_f7a9a92b[43]),
    .b(al_d6cb04b6[43]),
    .c(al_b8f391da),
    .o({al_98d4708b,al_5b8748c3[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_7241ba4 (
    .a(al_f7a9a92b[44]),
    .b(al_d6cb04b6[44]),
    .c(al_98d4708b),
    .o({al_e355574b,al_5b8748c3[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_f338b425 (
    .a(al_f7a9a92b[45]),
    .b(al_d6cb04b6[45]),
    .c(al_e355574b),
    .o({al_750642c9,al_5b8748c3[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ae399b3 (
    .a(al_f7a9a92b[46]),
    .b(al_d6cb04b6[46]),
    .c(al_750642c9),
    .o({al_ff2d726,al_5b8748c3[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_49e1e95d (
    .a(al_f7a9a92b[47]),
    .b(al_d6cb04b6[47]),
    .c(al_ff2d726),
    .o({al_53853e4b,al_5b8748c3[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_d5f8278c (
    .c(al_53853e4b),
    .o({open_n233,al_5b8748c3[9]}));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_b18ce391 (
    .a(al_d6cb04b6[66]),
    .b(al_d6cb04b6[67]),
    .c(al_d6cb04b6[68]),
    .d(al_d6cb04b6[69]),
    .e(al_d6cb04b6[70]),
    .f(al_5b8748c3[9]),
    .o(al_89b35cc7));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_df4e4f36 (
    .a(al_4bd1c0eb),
    .b(al_f7a9a92b[39]),
    .c(al_5b8748c3[0]),
    .o(al_3b7f0416[39]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_4c5ffe7c (
    .a(al_d6cb04b6[60]),
    .b(al_d6cb04b6[61]),
    .c(al_d6cb04b6[62]),
    .d(al_d6cb04b6[63]),
    .e(al_d6cb04b6[64]),
    .f(al_d6cb04b6[65]),
    .o(al_375b5a4d));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_1f5b6711 (
    .a(al_d6cb04b6[54]),
    .b(al_d6cb04b6[55]),
    .c(al_d6cb04b6[56]),
    .d(al_d6cb04b6[57]),
    .e(al_d6cb04b6[58]),
    .f(al_d6cb04b6[59]),
    .o(al_12dcd287));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_d3d9efcf (
    .a(al_d6cb04b6[48]),
    .b(al_d6cb04b6[49]),
    .c(al_d6cb04b6[50]),
    .d(al_d6cb04b6[51]),
    .e(al_d6cb04b6[52]),
    .f(al_d6cb04b6[53]),
    .o(al_ff1931b3));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_22c3e4e4 (
    .a(al_89b35cc7),
    .b(al_375b5a4d),
    .c(al_12dcd287),
    .d(al_ff1931b3),
    .o(al_4bd1c0eb));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_aff5fee0 (
    .a(al_4bd1c0eb),
    .b(al_f7a9a92b[40]),
    .c(al_5b8748c3[1]),
    .o(al_3b7f0416[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e71f9e45 (
    .a(al_4bd1c0eb),
    .b(al_f7a9a92b[41]),
    .c(al_5b8748c3[2]),
    .o(al_3b7f0416[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_1a3b62e (
    .a(al_4bd1c0eb),
    .b(al_f7a9a92b[42]),
    .c(al_5b8748c3[3]),
    .o(al_3b7f0416[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d0e883ca (
    .a(al_4bd1c0eb),
    .b(al_f7a9a92b[43]),
    .c(al_5b8748c3[4]),
    .o(al_3b7f0416[43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_4920adb7 (
    .a(al_4bd1c0eb),
    .b(al_f7a9a92b[44]),
    .c(al_5b8748c3[5]),
    .o(al_3b7f0416[44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3624d080 (
    .a(al_4bd1c0eb),
    .b(al_f7a9a92b[45]),
    .c(al_5b8748c3[6]),
    .o(al_3b7f0416[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_ee96519e (
    .a(al_4bd1c0eb),
    .b(al_f7a9a92b[46]),
    .c(al_5b8748c3[7]),
    .o(al_3b7f0416[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_6031dab6 (
    .a(al_4bd1c0eb),
    .b(al_f7a9a92b[47]),
    .c(al_5b8748c3[8]),
    .o(al_3b7f0416[47]));
  AL_DFF_X al_5fa3a508 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[0]));
  AL_DFF_X al_fed1cf92 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[9]));
  AL_DFF_X al_3e150ba3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[10]));
  AL_DFF_X al_b70fa3c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[11]));
  AL_DFF_X al_6feeb671 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[12]));
  AL_DFF_X al_c3966a3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[13]));
  AL_DFF_X al_65b28529 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[14]));
  AL_DFF_X al_e2654e41 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[15]));
  AL_DFF_X al_a72db636 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[16]));
  AL_DFF_X al_177c60fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[17]));
  AL_DFF_X al_b4d340d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[18]));
  AL_DFF_X al_e9eebab8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[1]));
  AL_DFF_X al_32ffbdca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[19]));
  AL_DFF_X al_3c74e279 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[20]));
  AL_DFF_X al_6b4e22ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[21]));
  AL_DFF_X al_682ef3b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[22]));
  AL_DFF_X al_8f5f4463 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[23]));
  AL_DFF_X al_b3eda49 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[24]));
  AL_DFF_X al_82e04 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[25]));
  AL_DFF_X al_2fdeb21a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[26]));
  AL_DFF_X al_41cbe38a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[27]));
  AL_DFF_X al_751ede8a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[28]));
  AL_DFF_X al_66bef662 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[2]));
  AL_DFF_X al_18f156cf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[29]));
  AL_DFF_X al_e19e0e17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[30]));
  AL_DFF_X al_b29d2972 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[31]));
  AL_DFF_X al_e34fa351 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[32]));
  AL_DFF_X al_19926c0f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[33]));
  AL_DFF_X al_5e4c14b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[34]));
  AL_DFF_X al_36c3eef0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[35]));
  AL_DFF_X al_fac75e46 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[36]));
  AL_DFF_X al_2c1e9112 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[37]));
  AL_DFF_X al_cd5f1797 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[38]));
  AL_DFF_X al_69a5c5fc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[3]));
  AL_DFF_X al_53439f4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[39]));
  AL_DFF_X al_11e6655d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[40]));
  AL_DFF_X al_13289cc7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[41]));
  AL_DFF_X al_4452d0a1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[42]));
  AL_DFF_X al_ed8ffd62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[43]));
  AL_DFF_X al_f6307fd7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[44]));
  AL_DFF_X al_e9523c4c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[45]));
  AL_DFF_X al_c8f61bef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[46]));
  AL_DFF_X al_b586de44 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3b7f0416[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[47]));
  AL_DFF_X al_1482b16b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[4]));
  AL_DFF_X al_171419ae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[5]));
  AL_DFF_X al_30889faf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[6]));
  AL_DFF_X al_aa222510 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[7]));
  AL_DFF_X al_68b359e9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_f7a9a92b[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_5283b07c[8]));
  AL_DFF_X al_79e10fbd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4bd1c0eb),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[0]));
  AL_DFF_X al_ed85ea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[1]));
  AL_DFF_X al_9470906d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[2]));
  AL_DFF_X al_7d9ad012 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[3]));
  AL_DFF_X al_ca41741f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[4]));
  AL_DFF_X al_e6a1aa76 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[5]));
  AL_DFF_X al_1a5b7218 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[6]));
  AL_DFF_X al_48daf472 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[7]));
  AL_DFF_X al_129c3e06 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_4dd3fb65[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_3cd0a9ea[8]));
  AL_DFF_X al_4aa179ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_36d845bb[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_4b6a4daa[0]));
  AL_DFF_X al_b6814fc1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[37]));
  AL_DFF_X al_ad8e28a2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[38]));
  AL_DFF_X al_b6e7e12e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[39]));
  AL_DFF_X al_798b7e68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[40]));
  AL_DFF_X al_c4599680 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[41]));
  AL_DFF_X al_9e476f67 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[42]));
  AL_DFF_X al_f1857961 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[43]));
  AL_DFF_X al_e7979d5e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[44]));
  AL_DFF_X al_df94c22f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[45]));
  AL_DFF_X al_1f65882d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[46]));
  AL_DFF_X al_f28df47d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[47]));
  AL_DFF_X al_88079c7b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[48]));
  AL_DFF_X al_a97be48f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[49]));
  AL_DFF_X al_29dd2b57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[50]));
  AL_DFF_X al_e5c54ba7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[51]));
  AL_DFF_X al_ab3b0fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[52]));
  AL_DFF_X al_8423475a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[53]));
  AL_DFF_X al_90b4c795 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[54]));
  AL_DFF_X al_1f170942 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[55]));
  AL_DFF_X al_f60ec6a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[56]));
  AL_DFF_X al_25e4d7ad (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[57]));
  AL_DFF_X al_fdb1f1c2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[58]));
  AL_DFF_X al_645997a0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[59]));
  AL_DFF_X al_c069c7f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[60]));
  AL_DFF_X al_aef45de5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[61]));
  AL_DFF_X al_758ecfdd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[62]));
  AL_DFF_X al_4e73e7f0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[64]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[63]));
  AL_DFF_X al_ddb6e4d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[65]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[64]));
  AL_DFF_X al_a9e6ca42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[66]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[65]));
  AL_DFF_X al_64bc980d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[67]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[66]));
  AL_DFF_X al_b00817e2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[68]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[67]));
  AL_DFF_X al_588b0fb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_c1960abd[69]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_6f9059d1[68]));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    al_c9b54fe4 (
    .a(1'b0),
    .o({al_ac55c9d9,open_n236}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_fcc311f3 (
    .a(al_5283b07c[38]),
    .b(al_c1960abd[38]),
    .c(al_ac55c9d9),
    .o({al_869b4e37,al_93772c3[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_2e616347 (
    .a(al_5283b07c[39]),
    .b(al_c1960abd[39]),
    .c(al_869b4e37),
    .o({al_ca5ea173,al_93772c3[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_dfd6cd89 (
    .a(al_5283b07c[40]),
    .b(al_c1960abd[40]),
    .c(al_ca5ea173),
    .o({al_76985513,al_93772c3[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_58b1fe20 (
    .a(al_5283b07c[41]),
    .b(al_c1960abd[41]),
    .c(al_76985513),
    .o({al_8b8db5a8,al_93772c3[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_53aed3f9 (
    .a(al_5283b07c[42]),
    .b(al_c1960abd[42]),
    .c(al_8b8db5a8),
    .o({al_8d3dc6f8,al_93772c3[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_9fc41504 (
    .a(al_5283b07c[43]),
    .b(al_c1960abd[43]),
    .c(al_8d3dc6f8),
    .o({al_af8cdc32,al_93772c3[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_14fec680 (
    .a(al_5283b07c[44]),
    .b(al_c1960abd[44]),
    .c(al_af8cdc32),
    .o({al_50432123,al_93772c3[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_ddb1f0c6 (
    .a(al_5283b07c[45]),
    .b(al_c1960abd[45]),
    .c(al_50432123),
    .o({al_2637e6b1,al_93772c3[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_4492554 (
    .a(al_5283b07c[46]),
    .b(al_c1960abd[46]),
    .c(al_2637e6b1),
    .o({al_d2ba203e,al_93772c3[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_771ce68d (
    .a(al_5283b07c[47]),
    .b(al_c1960abd[47]),
    .c(al_d2ba203e),
    .o({al_72aa54c,al_93772c3[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    al_bb4a8d29 (
    .c(al_72aa54c),
    .o({open_n239,al_93772c3[10]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c8b4744b (
    .a(al_8b60a1f7),
    .b(al_5283b07c[38]),
    .c(al_93772c3[0]),
    .o(al_bcaebe78[38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_d2db202d (
    .a(al_8b60a1f7),
    .b(al_5283b07c[39]),
    .c(al_93772c3[1]),
    .o(al_bcaebe78[39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_7d85a6a0 (
    .a(al_8b60a1f7),
    .b(al_5283b07c[40]),
    .c(al_93772c3[2]),
    .o(al_bcaebe78[40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_cb483c2 (
    .a(al_8b60a1f7),
    .b(al_5283b07c[41]),
    .c(al_93772c3[3]),
    .o(al_bcaebe78[41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_79bf8fd7 (
    .a(al_8b60a1f7),
    .b(al_5283b07c[42]),
    .c(al_93772c3[4]),
    .o(al_bcaebe78[42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_e81a4d38 (
    .a(al_8b60a1f7),
    .b(al_5283b07c[43]),
    .c(al_93772c3[5]),
    .o(al_bcaebe78[43]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_63354f7f (
    .a(al_c1960abd[64]),
    .b(al_c1960abd[65]),
    .c(al_c1960abd[66]),
    .d(al_c1960abd[67]),
    .e(al_c1960abd[68]),
    .f(al_c1960abd[69]),
    .o(al_5c60fab));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_186b4c4b (
    .a(al_8b60a1f7),
    .b(al_5283b07c[44]),
    .c(al_93772c3[6]),
    .o(al_bcaebe78[44]));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_f461cf7 (
    .a(al_c1960abd[58]),
    .b(al_c1960abd[59]),
    .c(al_c1960abd[60]),
    .d(al_c1960abd[61]),
    .e(al_c1960abd[62]),
    .f(al_c1960abd[63]),
    .o(al_aa0aca8a));
  AL_MAP_LUT6 #(
    .EQN("(~F*~E*~D*~C*~B*~A)"),
    .INIT(64'h0000000000000001))
    al_68644f10 (
    .a(al_c1960abd[52]),
    .b(al_c1960abd[53]),
    .c(al_c1960abd[54]),
    .d(al_c1960abd[55]),
    .e(al_c1960abd[56]),
    .f(al_c1960abd[57]),
    .o(al_26b3b41e));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    al_b65ed13 (
    .a(al_c1960abd[48]),
    .b(al_c1960abd[49]),
    .c(al_c1960abd[50]),
    .d(al_c1960abd[51]),
    .e(al_93772c3[10]),
    .o(al_27f44dd8));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    al_61cfbabc (
    .a(al_5c60fab),
    .b(al_aa0aca8a),
    .c(al_26b3b41e),
    .d(al_27f44dd8),
    .o(al_8b60a1f7));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_5d17b43 (
    .a(al_8b60a1f7),
    .b(al_5283b07c[45]),
    .c(al_93772c3[7]),
    .o(al_bcaebe78[45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_c5f3e6d2 (
    .a(al_8b60a1f7),
    .b(al_5283b07c[46]),
    .c(al_93772c3[8]),
    .o(al_bcaebe78[46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    al_3f7a20f1 (
    .a(al_8b60a1f7),
    .b(al_5283b07c[47]),
    .c(al_93772c3[9]),
    .o(al_bcaebe78[47]));
  AL_DFF_X al_7bcf5218 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[0]));
  AL_DFF_X al_210a05ef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[9]));
  AL_DFF_X al_cd8e639f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[10]));
  AL_DFF_X al_7ee8e1ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[11]));
  AL_DFF_X al_185c12f4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[12]));
  AL_DFF_X al_b6cf0894 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[13]));
  AL_DFF_X al_4f49e6be (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[14]));
  AL_DFF_X al_2eb20435 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[15]));
  AL_DFF_X al_1321fd4d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[16]));
  AL_DFF_X al_de1fd319 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[17]));
  AL_DFF_X al_b21eb769 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[18]));
  AL_DFF_X al_567a7cda (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[1]));
  AL_DFF_X al_7b8950c7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[19]));
  AL_DFF_X al_a7666c57 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[20]));
  AL_DFF_X al_85d2e651 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[21]));
  AL_DFF_X al_1f1de636 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[22]));
  AL_DFF_X al_1fecf4a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[23]));
  AL_DFF_X al_af217015 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[24]));
  AL_DFF_X al_a05487f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[25]));
  AL_DFF_X al_359627aa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[26]));
  AL_DFF_X al_eef974cc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[27]));
  AL_DFF_X al_91ce5b89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[28]));
  AL_DFF_X al_4ed4b91f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[2]));
  AL_DFF_X al_2fd4cb65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[29]));
  AL_DFF_X al_dcecf5eb (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[30]));
  AL_DFF_X al_6b5e0cae (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[31]));
  AL_DFF_X al_348599a7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[32]));
  AL_DFF_X al_c5d00881 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[33]));
  AL_DFF_X al_7914ac65 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[34]));
  AL_DFF_X al_863c752c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[35]));
  AL_DFF_X al_b87671ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[36]));
  AL_DFF_X al_3a84fac7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[37]));
  AL_DFF_X al_1b6e7fef (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[38]));
  AL_DFF_X al_3ba6d592 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[3]));
  AL_DFF_X al_528c69b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[39]));
  AL_DFF_X al_91bca1b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[40]));
  AL_DFF_X al_d8b3ca1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[41]));
  AL_DFF_X al_de95278d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[42]));
  AL_DFF_X al_98f90e2f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[43]));
  AL_DFF_X al_314cd44c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[44]));
  AL_DFF_X al_74c99470 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[45]));
  AL_DFF_X al_c2ac6352 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[46]));
  AL_DFF_X al_8abb52f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_bcaebe78[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[47]));
  AL_DFF_X al_80a6f628 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[4]));
  AL_DFF_X al_e1d4e1a5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[5]));
  AL_DFF_X al_a685201f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[6]));
  AL_DFF_X al_9b6cdee4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[7]));
  AL_DFF_X al_d4982e74 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_5283b07c[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_f2b51288[8]));
  AL_DFF_X al_a32a67ca (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_8b60a1f7),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[0]));
  AL_DFF_X al_7bb68e0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[9]));
  AL_DFF_X al_67c11257 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[1]));
  AL_DFF_X al_79808e2c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[2]));
  AL_DFF_X al_96dad4d3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[3]));
  AL_DFF_X al_a6c245fa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[4]));
  AL_DFF_X al_1fab1a62 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[5]));
  AL_DFF_X al_4d31daa (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[6]));
  AL_DFF_X al_41689714 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[7]));
  AL_DFF_X al_a324b997 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(al_3cd0a9ea[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_fac191b8[8]));
  AL_DFF_X al_69b4fe12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[47]));
  AL_DFF_X al_47547ec8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[48]));
  AL_DFF_X al_673c5a1c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[49]));
  AL_DFF_X al_dd16212d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[50]));
  AL_DFF_X al_d824ff53 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[51]));
  AL_DFF_X al_80f6610c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[52]));
  AL_DFF_X al_323be77e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[53]));
  AL_DFF_X al_80dc8452 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[54]));
  AL_DFF_X al_3661ca68 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[55]));
  AL_DFF_X al_fecd4530 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[56]));
  AL_DFF_X al_458d9ab9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[57]));
  AL_DFF_X al_937eff72 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[58]));
  AL_DFF_X al_d751125c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[59]));
  AL_DFF_X al_23bcfb1a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[60]));
  AL_DFF_X al_cf76943e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[61]));
  AL_DFF_X al_1d68e107 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[62]));
  AL_DFF_X al_7157cdaf (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[63]));
  AL_DFF_X al_70a1b090 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[64]));
  AL_DFF_X al_d7efe57e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[65]));
  AL_DFF_X al_592eb0d6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[66]));
  AL_DFF_X al_9d5a1699 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[67]));
  AL_DFF_X al_de9867e6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[68]));
  AL_DFF_X al_d6194c5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[69]));
  AL_DFF_X al_4f71f3d8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[70]));
  AL_DFF_X al_bdd30786 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[71]));
  AL_DFF_X al_76df1b58 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[72]));
  AL_DFF_X al_f420246e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[73]));
  AL_DFF_X al_a28f682 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[74]));
  AL_DFF_X al_6e8db4fe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[75]));
  AL_DFF_X al_47dfd70 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[76]));
  AL_DFF_X al_1870bb89 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[77]));
  AL_DFF_X al_c156871a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(denominator[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_9d1d5c0[78]));
  AL_DFF_X al_35b11324 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_dc871c53[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(done));
  AL_DFF_X al_bb2a0a10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[0]));
  AL_DFF_X al_c3812f56 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[9]));
  AL_DFF_X al_686f20db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[10]));
  AL_DFF_X al_fcfebea6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[11]));
  AL_DFF_X al_7732f4ec (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[12]));
  AL_DFF_X al_f3f58b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[13]));
  AL_DFF_X al_e61c4c93 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[14]));
  AL_DFF_X al_6a73ad4b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[15]));
  AL_DFF_X al_1ac47d42 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[16]));
  AL_DFF_X al_3e9294ac (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[17]));
  AL_DFF_X al_5668b702 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[18]));
  AL_DFF_X al_75b89d0e (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[1]));
  AL_DFF_X al_cd57881c (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[19]));
  AL_DFF_X al_9506411b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[20]));
  AL_DFF_X al_fd541c99 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[21]));
  AL_DFF_X al_9e70e012 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[22]));
  AL_DFF_X al_5b158070 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[23]));
  AL_DFF_X al_693bc92f (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[24]));
  AL_DFF_X al_e7396a48 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[25]));
  AL_DFF_X al_3af3f245 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[26]));
  AL_DFF_X al_708041c0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[27]));
  AL_DFF_X al_bbfa7acd (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[28]));
  AL_DFF_X al_1d89aa25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[2]));
  AL_DFF_X al_eba09a4a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[29]));
  AL_DFF_X al_7e47ad43 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[30]));
  AL_DFF_X al_f30d22f6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[31]));
  AL_DFF_X al_377a57dc (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[32]));
  AL_DFF_X al_9737e66b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[33]));
  AL_DFF_X al_bc8da1a8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[34]));
  AL_DFF_X al_67350fb9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[35]));
  AL_DFF_X al_3652fa83 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[36]));
  AL_DFF_X al_35f523e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[37]));
  AL_DFF_X al_fc6db617 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[38]));
  AL_DFF_X al_bfcb957b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[3]));
  AL_DFF_X al_929077a (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[39]));
  AL_DFF_X al_41a25649 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[40]));
  AL_DFF_X al_9da157db (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[41]));
  AL_DFF_X al_d3c7356d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[42]));
  AL_DFF_X al_f5583890 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[43]));
  AL_DFF_X al_7741cd5b (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[44]));
  AL_DFF_X al_469fb578 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[45]));
  AL_DFF_X al_d1a308e0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[46]));
  AL_DFF_X al_2ce98575 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[47]));
  AL_DFF_X al_f3d4028d (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[4]));
  AL_DFF_X al_a6dd3266 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[5]));
  AL_DFF_X al_75f33271 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[6]));
  AL_DFF_X al_8c7a1c1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[7]));
  AL_DFF_X al_8140f785 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(numerator[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_a5806bc7[8]));
  AL_DFF_X al_211928d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[0]));
  AL_DFF_X al_a875d850 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[9]));
  AL_DFF_X al_b59bb075 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[10]));
  AL_DFF_X al_1a2500e5 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[11]));
  AL_DFF_X al_42bc6562 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[12]));
  AL_DFF_X al_ac4b7df6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[13]));
  AL_DFF_X al_71242670 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[14]));
  AL_DFF_X al_b3f0dfb6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[15]));
  AL_DFF_X al_c3ea0bbb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[16]));
  AL_DFF_X al_e44e8a84 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[17]));
  AL_DFF_X al_96a4b8ba (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[18]));
  AL_DFF_X al_46a2af83 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[1]));
  AL_DFF_X al_88f0f9e2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[19]));
  AL_DFF_X al_667462ac (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[20]));
  AL_DFF_X al_66b8286f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[21]));
  AL_DFF_X al_9b3545ca (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[22]));
  AL_DFF_X al_a8aa46e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[23]));
  AL_DFF_X al_fb14e4c6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[24]));
  AL_DFF_X al_c049dba0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[25]));
  AL_DFF_X al_4c960124 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[26]));
  AL_DFF_X al_a883ea3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[27]));
  AL_DFF_X al_c4fa88d2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[28]));
  AL_DFF_X al_d42e6219 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[2]));
  AL_DFF_X al_dbea5ac2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[29]));
  AL_DFF_X al_7c806850 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[30]));
  AL_DFF_X al_7af3ba3e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[31]));
  AL_DFF_X al_90b512 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[32]));
  AL_DFF_X al_6db674a2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[33]));
  AL_DFF_X al_58cddbec (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[34]));
  AL_DFF_X al_cc282882 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[35]));
  AL_DFF_X al_e7dc5b56 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[36]));
  AL_DFF_X al_3a805102 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[37]));
  AL_DFF_X al_3a0f8181 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[38]));
  AL_DFF_X al_4dada817 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[3]));
  AL_DFF_X al_f49a7269 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[39]));
  AL_DFF_X al_ff0133ce (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[40]));
  AL_DFF_X al_769dacc6 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[41]));
  AL_DFF_X al_903748b4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[42]));
  AL_DFF_X al_fb6ceb83 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[43]));
  AL_DFF_X al_df8911cf (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[44]));
  AL_DFF_X al_430d0ba1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[45]));
  AL_DFF_X al_a0b2215d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[46]));
  AL_DFF_X al_2c8dd00 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[47]));
  AL_DFF_X al_c3679cc8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[4]));
  AL_DFF_X al_67e73dee (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[5]));
  AL_DFF_X al_60987264 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[6]));
  AL_DFF_X al_a632a9cd (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[7]));
  AL_DFF_X al_87e3c4ed (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_3b63a678[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(quotient[8]));
  AL_DFF_X al_5e3d5ef (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[0]));
  AL_DFF_X al_53989262 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[9]));
  AL_DFF_X al_ec8df0cb (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[10]));
  AL_DFF_X al_cf9ee80f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[11]));
  AL_DFF_X al_307971a4 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[12]));
  AL_DFF_X al_1dc36712 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[13]));
  AL_DFF_X al_ad56177e (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[14]));
  AL_DFF_X al_c925149f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[15]));
  AL_DFF_X al_c39c015c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[16]));
  AL_DFF_X al_4f2f24c3 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[17]));
  AL_DFF_X al_d4f5a330 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[18]));
  AL_DFF_X al_4ca2f6e2 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[1]));
  AL_DFF_X al_73dbf462 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[19]));
  AL_DFF_X al_fbc71faa (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[20]));
  AL_DFF_X al_b074c41a (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[21]));
  AL_DFF_X al_d3914004 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[22]));
  AL_DFF_X al_e88f4dba (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[23]));
  AL_DFF_X al_1bd9f325 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[24]));
  AL_DFF_X al_132e504c (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[25]));
  AL_DFF_X al_b3f008f1 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[26]));
  AL_DFF_X al_794ced (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[27]));
  AL_DFF_X al_959fef33 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[28]));
  AL_DFF_X al_a7e80b5d (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[2]));
  AL_DFF_X al_f831e8ca (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[29]));
  AL_DFF_X al_890566ee (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[30]));
  AL_DFF_X al_1d45ea0 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[31]));
  AL_DFF_X al_c3cf0fae (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[3]));
  AL_DFF_X al_c107bff (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[4]));
  AL_DFF_X al_7e423429 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[5]));
  AL_DFF_X al_ba2474a8 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[6]));
  AL_DFF_X al_4ba4e538 (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[7]));
  AL_DFF_X al_fc2e9e8f (
    .ar(rst),
    .as(1'b0),
    .clk(clk),
    .d(al_bfaf4e7[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(remainder[8]));
  AL_DFF_X al_f6de6753 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk),
    .d(start),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(al_51794c84));

endmodule 

