


module mipi_dphy_rx_ph1a_mipiio_wrapper #(
    parameter LANE_NUM = 4,
    parameter BYTE_NUM = 1
    )(
    input wire                             I_lp_clk,
    input wire                             I_rst,

    input wire[8:0]                        I_clk_lane_in_delay,
    input wire[8:0]                        I_data_lane0_in_delay,
    input wire[8:0]                        I_data_lane1_in_delay,
    input wire[8:0]                        I_data_lane2_in_delay,
    input wire[8:0]                        I_data_lane3_in_delay,

    input wire[LANE_NUM-1 : 0]             I_lane_invert,

    output wire                            O_hs_rx_clk,
    output wire                            O_hs_rx_valid,
    output wire[LANE_NUM*BYTE_NUM*8-1 : 0] O_hs_rx_data,

    output wire                            O_lp_rx_lane0_p,
    output wire                            O_lp_rx_lane0_n,

    input wire                             I_lp_tx_en,
    input wire                             I_lp_tx_lane0_p,
    input wire                             I_lp_tx_lane0_n,

    output wire[LANE_NUM-1 : 0]            O_lane_error
);


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
jIH9ZrLe/lM0mD4RX4uCeQlIRk/gaZ9c9YFj8J2vJWtqs8Oab0xHT0t5lQin9jS0
QALf1v4RWPLqNQ1PaPozxPrr5r8Yx5kWJUVIAR0SZW0Fr4J1vD2UtsYrmzrr4qAE
0rFWsnDf+TQ0rTz96k+Ga+TDCnrKaVaWoySj1KsnFvA=
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
jGi0TY44lEethqDNUJvlgvGg//HrJEJCumcU0F+57ZmTYgEBHPqfOeJWBVstT3uj
oG28CF2PnxEENhFtgxpW2MCs4L5NM2Y19wAtUXazX1DPtIqSo1sgXdmzSLD3ce+4
dRACUBJKPrd+TVn4cvZkW2N5OyV+9pFSo4Xqkcpa0vo8l9uETwwARC7oBu0v4ngF
QE7ExxGWDQqjgZCUyz7BB54w5/gMuGIpLcY+LVfXdmu+DJ5chFs0tdukrG7rXx14
0QBe4W2hv8rKtKY6O2HqApCvxjGEZ5UhJAK1Xbu5kABTYfhSnJSK7iTlEyiFjCqc
efmYTicyeStQ4a+9sjYtWw==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
AgiXzKAt0yDAatE857meJJRn0riDoGEnOnA2wKJIrW7x6Rmx1RBQgR0pRARCiv4Z
d/JsOEpZIQ8HPlvO9O7/v9ybsBJRWjbeS2xBFJyW9ZETdp8qg46sT+8mJYeJL53M
JYRDMf/Jn8on2yFDC1MhdI0YZpmHp6241WTnpdROyZQ=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
D5SfoLWugiUy6Nh000SkkyZr+2dqCGFclh+5SNINQkVu5bcDCUM3i3seD75v1hFl
/9XCipLqiMEkiP7KxnhQN5WtaCHLBBAMVNRayhbTbu9xtR0F6H6/YhRsfwkiibMZ
OFQfUJ+ECqVEu7mUQHCw4X5CwQxpf0ZkPsvUk3t+WrCDFJCy+QWA4anQq4LTnpwm
yUffXifqu2nd6pQjayhtFWUT68O42LyqeJYRNfP8/mihHsvVdCY99q0npGJNZ6y2
zoPaGDyYfIrzlUJs7gfTduPQMW8LJm0VqXS7qiaTX5AR8+Uj3CpBb4FehpcyA1x7
G46thGYGcdSMhiFZE/dKNw==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
jQrBJ/bJXCnlMyCNXGJOwYYWkBCOzCYKJqKCCWFtqvrAbcWzpyZ3gYqLt5E471uL
TZhkpwBHTFJQ+tnhrGIF0pddW2drzczv9TEVgUVMw5VYp+nazsH5zEIxUbhlvGmM
lAsl/EO+E4Lcwg91aN3ULer3dIULdw1soCCAEMcg7Bw=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 43216)
`pragma protect data_block
vP0bRwUKZ31KeD8aAWZKClJYNPg1a36sVVcHoej6aT6MP6J0v0m3K6Q2L12o661E
sMySLpeqLN6vj2dswxMWY1MmPDQg7/lVr78wDGzm/JfHl4ec2hw0C/Je0LgGvnWJ
442+KJfBFFvjDvSN3kUz6mYD/2F6iV3o9kCx5fvWprS+0VT6pe6gU0/1b7VDZ/nV
6mnvL0qKNMuOL4Y5slnKF/f40l6Z0W0jjBXf+ZpOolSloaVJMhXbJuevSB+a6KoA
Z/Z91/7Afb5RmzSLUjkmR1zeiq2Ew4oESqjEQIXtzh+tf68st2TbM5fMbwx6D5z/
LGEIPFzuUrxPFckytHolC/rPM+RcnpGEgH5MF2S0HKoQUBkO2D3FDh+0eiZBP/OO
HDdp3duucIG04Y8at04f/mearLbFgI6AvN3XbYl4mSU8irb/c6AgGcK/mgUUUBDK
khz+S3Zj9Kai4l4kvmJvM9cNcF9j9zKqsSGDTtfLUgaNB9B/GulieGHm5lZec5xy
TQWhyyPGQPtc2mJQlY59wR6ZYuUrZxg6nQzTSP2IvjKzkfzGDSioqsolH1iYHAxm
iu8WczDKN9LQCXprmb9bKCCug/iSQB4y67/CYSBWaO7g1cv9hKYGawZVGumWHvxM
aQK1kyx1Y9bV6gTMYHXixqkh/Fpa/0ik5zuRNZbxeDULxNc2iTce+yTeJwvE0lfg
uZujDeyfzLyLTFmp4HAUsISaewhnfhFw+J3TKMFDFkA91ruDAvIOq3SUC3x80ng1
aCov4d5chdHfGsmxwbF0Yw4IIa7p5qFupM6bW71bkFw75VhiPfWpdGF2ED9ydJrI
WxBvibijzIvjSrpzRaP5GM7ewNpAFLIaWUc8EpKcePk9ZtqiHn37reIoJTnc3dbk
EQJZYKOrMrSpMm7nIc2Jbh4BNpEgjyYTC9Id07PEqjxr8tu1MaN4py8Ab1r5386z
GW0kBVxFwGkmSXfzgdRa6c0awUEPp5dO8gmKSZDo4XB3n2PwMGdnthFbK7jCtDUm
62U425E26kUjOrTuqf9IOlHQt6P7QdEKt7mF9VvB+x2wn4YRmMLlCUGcMSXy5U+7
Rn8adDBMz85ytfOsL8I1oomv/0rxKdRXiPNaZFLghQtyq5REffTHPY893HUUO5eZ
gBQt4b3kDEZHxyK49mxah5Qo+uCEbn7lztsQDN56X6frhYVTko3VoVHmYxqTgM9D
V6ZFFd2ntmkYulGBcT4TU+ojMQxzlk154FCOcN4Fu5ynFoR0v8HHg5h3XFKHZwWV
Y7c9SoYlljQew8j34qpKSAjCNCtOUZSKIlFWhkYIJ6ERDg8L+75EHwZzVU3NCWuh
1GZode2O7eQ1aAdKmrdmX3O4CUwcOF5UgwSkw2U44oEeCl12Y7Ar/Qp+/ar2SJ5/
o/yjmiVLpVHOt2r7EaqiFD6UUZ0c/gaHA5NTDgWeTBMDHQaslecDwb2rN65MVDV5
Ia3Tl+EfrPWZ/oggycE5r0I86Bh04n17DzKflGQvT4axY047PbTgpe+qaFg+aCKE
nB2Ky8QjZQKQ6zgYidZyrAkFcfy+8Gik3paA4OaT2sU9pzDaf1iwewdyNpyq1NXs
5/9pZHbpa9+jbDNLIaidBfGuQReTTMQKoWOdl2hoIVckgPeXgSwMbvMm/AReNT4E
P2sqHQ2aAeq6Y289AQS6CXHnEQOUjdT7dwAOe/6z0AvgZGDV9WBAncYBaxR1E0zE
rhScb4wVr/RS3SKE18nFKk347nVMgE8p+gMJVtCGqclzj58rHqyqH6S3sEwG0d66
eTwkMpoc1yrZbouIJeiD7141suV8NDjHVtrAM6bPqVWpWai/d3cqzzxXm6t4jHcI
KF1p1rhdbz6VlArbQR2O9fq270fQrmfLiD9wtPtcZQRHI5yT7wLBkNKOlerK27co
lYbmi91GkQi/nn4YB0t5oHAU0VnIrrv1nZZHstX3Rh51sol4J/+MfJpSLAJxZgp+
Y2hUOn0iCWXMlNL93IZ8kbjosZyIcdFo6Gv6+Cz7HaSkerDjwqPo3adkRlnXZ8J0
Pau4+W+6xGSMipizaZUbVMjzB/FLcMrEVMD71CgUWh1pedOIdTx7hIOMbFWupdyt
JnHOLppW7e1Is9A8bcfWDgBc33TIvF6PzV2yBEM9cOPvGXwbzGMG+vsiOaTRVsF0
roOv6dccH8bOv8oBcCPkRRWBkSki0Z66jeJaEUx5eFOq3gKgBDUxe7g5tcSLnMLj
Fw94r2qklgELltw/Ew3AaqEjiPjZUb6LF33VinOMVD3CgT/vzHBN7Llw3SUD6xIP
lhr1NV15aO6e2nhUy4orO8AcX8NGJr6WH2R2xFU3DPKdaiZJZbCdn/EgFr5MczyG
QTAgdBSk0UoZMB0n2KDXLQOaobZaD0nkIBcctIyAzbO9sz3ts0DJk47x6He7wk5W
CRVQTBQk5DUHVvDyfady4/36QoRM2YUYdnFQ7IZ3VX0bitY+pmH63Xiy2ReWM+Sw
eKajNVKkuz751VRDOa2UbXLyF/LxaaiXs+064EKxbBRIpIHAhuttX5XHD7EIs0VJ
O4+6kWulU6cUVpleevGlp50U7ISKi6AYuT6vaWyUYbmElLpRUslGeNiJ80SOe7uL
I1fIwwtoD9eZ6wFEDdpd8r0G08PpVcNvzxnAXRsdGMu3WgonoNiixBID7eEk51hf
DNNICHOBV41r4zn3Ud2NlBkzxWeDO2OkzTQjvXt9o1nRcxfwdI8pfSf5O2bgdLqS
d2Uji1KjgIRrsqtTpjOJgiCkdwOrC2S1puvjA3d7gd85DS5pAFqpMaxjBibmpSCP
yHQ1I/JQJIsxZLD0sAan6f5LLZbu3zvJgi6DxJy4kGgc1uF1WNBOknlUn0EJPP8t
1qnICGES7yqVTrpY7/NnYvannQFt+GA+XtSnr4D6JfRrI+6Bepm2JTiVebesOKzd
8ChKC0ewVderwGi898ZGvnQfcCSYcMjcL9eGbQAj45WfJK5R20qQob1wVtb4cSId
35iWGVwJ94jwg+EeufNgeQP1sq1ABlulXemlNV1ungV5SY82po8Omkt4/xLU1CrQ
OVtIr7CMvo4WnIZiua9YQEHwvqtPIOOyvzrfgYHmTiromalanFZWmMNC01wlMzgj
mxCIvV5srCp32MeNdiOaOeSxCGF1ay0kw14ixrHkjZUrfjYhhj6wkk2WiIy5RDj3
3ScEH5rCoa3bwMpxC7qd9tnCi79GmUDLlGsMdopG0agG7/361fhy3I4x2pWY4TA7
4d8aymlBr1kXIGYm60IHAvy70N8PxxcjvXbOJvLKjBygfH7zzNvOVOiP7HFH3G/p
+g3cgmOl61PhnndrlYyyr9gl+gy0cKjUoJDI7m/73tomoBAwwRBJ4h4miXmwTHg4
dK4i1ugx6gQcGCBSJJ13SEKA+M7scDksCl4VZaL/TiaqqR3dQFsiWJYmRmoF0GXm
dPiz5h9Lh9ENyygV2/Gn7a55GmHC+nOimgegBywZYiwqbDIi0lfZK09aYTpFDSBY
v6FPleZJwW9kFe37qda+0NcFB+TsDCS89/xEdc2Fd4tRogbQb6ow0XBb3FW2OrU3
u/qEaE90RFfYyFtSh6DPw5P81Yn1NDjVg3iNp13zEkcOfcxADOfacS8uZlYePU8L
oQTsX9lGXTWL8kOXRclEdwfArmcFbzQ0ZsoXnFSwohpJsotux9hl7l23KWTB9f0G
4pnA27sAlIGAjVri5x7hoocLen6LZd/HFpXk8EFBlAKquSCmoAfP9YDz+IqGmAwA
eDPa1CJ/0s1Y3LLlW3eLZGwoa9lkfpmzax9n+IcME2oRChHeMi/f+tsj0LAbHgIi
GpW14MV/5Hc2WiaOBj/4uhx7Socv4rr6zRLe4+Np4hVWyJyw5YZIjYTm7KN/I5AT
VqaU0+JdRO/fcfNmSNKYo5Y0kiieXq/tLh7++fSanhhu5nAQcUG6+xOt8ze14oJ2
Cl7u9lINXgPNh35CDb5LSbgSRAPlx5EV2nZUnAyudj17kZdQKRFpviWdYIZbSxY6
kIuxYlA08mwkwCf3QKSx7thOV2DMjELVh2YujfUE596xp0QKhotO1pLELJg/MWTg
qPjWyQ3ePQQWfiFyRKDeXmDg2DhH0kHIARh2V56n4bW+Z8mx1e2oPMso/qqr7Wpo
iypqE/VrqLGXYC2FC+L8HyICa0t0Gxu4kNT2JvhE9f2m37mZC+3+dc302vm+7XiT
/aK8A3EyEtH5CnwyHDHbhxlEHnB86iphpO+FEFqeOFpJv6Oz+pYU+/YFBnV3z2D3
gtfXb4L+gu5Jc5tetKcKmqluHVwL/NrPpf2AWCJwuw8/oT0rrw6WYua8yHzEmXHv
6BuvVZthUv7s71VQ7EsVEVXOsue/ktrPeXFSzkwGewsjKx5QPGbSbU/2588j2nYn
wwmoczO602j8iBvuijm5z8LmzjZFSvM89w+gKbkLVDaxGKhNHAqUJ09i7zsg3fHb
BAytvxN5bria7r6D4TMxnJDGDNGtVzFqalyIgrZlVbmWfSloM9SvuyJYX87QV8Wr
FWYZq9PKBaMejJRwDxrtqmMXB3gpwc49jk2jRb8PKE7hp8Oqt5+UOTs+RCdNZlJ6
O/CVHgYJuhVh5c0OUC29kJV74cRb53Oe/XL0ZexmgIX+pwd0GNy01XlxqH+oeLT5
lf7gOHz/IyCclUEs52se0qXOj7g6FZmQ0kvu0NlZMY6Vz7yoXDnpV6gim8YrOIOd
zgYwpdzmKS9Bw9dyryFem6wHSn6M/7RODGfu+ARpRRvQNZt81aduiCboI+qH5CEi
VVMKpieFmb/TtOMDRWq+7tQ11rTiuENJ8ZmVPsYLAvZ6MhcWzT1u/hRHwh2m68rn
eId8Mz8V4L1zzXb6ZwC73xbAlpqxn8gcXond/o448vR7C44p6ux4OkmHavf0Av7r
XMAxQfAXDabPlyANlp8cHYY9LmNOeH2SI+DGj6DkstW4Amd7sCAsv1Y0LdQa177Z
ql1PyxlOgck841YVPZFp5DhFkROWF/Ysc82sd50SndkjM1G8exFhxBFEXhV+5dA/
km2+DfylQVbOc2xxwFlPTLxmbkwicZx94Vgp/eXLJ1kx4Ngh0AEA0ODImx5OWsbX
mk8DlCZbvwNaxT9N7m9++EQh+z6enFMolzbHPV6SE5QEaWByfdlAUoL5zXG2SxoR
gp2OQsFQtGfge5cMrha/K6G8v3jC/v3uG1VyZQDvfRWeVr3uNg8wVQm1y9TrCSq0
+ZT4foKK0TlygEgOaoIKk/bIMmrvAKQhXY2KwEawSNXC6Q2Ca2AH7c3Qu6oFVQgU
Z4wRIak0XjcMgOpxO/wFPaZQVhiRvt8bJzG9g+uRPdaTytbiXSrcz6frtbBOmHGs
SJRoCSH/Gl+/JlmyS8SXcBNWTv63l185hpGq8QaDLe7NRLsfsfWkZjcC5wrHSyPJ
oMQxR9PppOiYKbAqIk3hSc3XoXYipD3GuGNN7qBXQmjy0UR2+MXAojOD+T4w1asQ
lGSBRi/YVMzmyp2BqPkMGJ8uoDqYeyReRmkaMFaM/0dhylWgdGMdvq5gclCDUIR7
Z1HGTbxwwPLzVAks6TRVKdJD7KsCzQ3iVlCjErhMrfJAO9mVtpCtVipzYfIp+qLq
txslWqFAKQWvSlrgwphwsO9Oatxy/f56z8ScD3jXPrA/9XQdiPk+nO05frNgyebm
netkWeTcgaY2N1vfj9ogtVKOWKyA5rOcU+effJuWNfLCQBhCVlZawix0uKDAXCdw
+yt1fbFOF86x+ugBl8mhyiR8irvm7H7Wt+I46MiaYGI5jXmgZ8Dxqu4Ggy0KAsT4
PwP2d9syq5NUNz1NcY0ZhOR1Zn0C/2QMN7uWOqXyFjnjidB5gD0jhv2VnWKIVlGX
GmMyK2hfoG60jOBdP9tcHIeMigF3+VpANiKyVftdc42+Qpg2r9BRGPMZ9gjJHycU
ng11+MEGT8hltLTY24eTisNvquwqDztPPg8qDrPDKDNdpsdM8fGx74xx1q940V6Q
T3xVKPkIZsAbfLB8TpGavjakTEo8xlUTlX078p+cuyBaNZ0c7+7DsXO7+NnZgOX1
O7xzu2AXuZmODoicawDi+wHcrvn2mPKubV3qR00FDIeK1mpheWw13D89w8uVKnXP
zdh3fQZIG7r7Lkb/vtoH8AYVEHa1iVCknPXTyL3DuZtFJvYuxwQFxxemr3sWqN4l
f+gawCeh7zsqD/qNa0OSt4osu7X7tP6L/vmXjf39dyXcdytKlvEKcHgEMCLf/Gtt
sivaSyzO4VYgu8fU6ytAS+OYKikAtOcy1yijQRF5LZyfERZ05FT0OiZKJ0CKjc9W
XH6on5af4IFkTySUWrHu4XYI0/sQnuN7ZPOqo+xht/nGsQ6kf0qOLuhRVnjx45Nw
G29SERm1DL6S1H2deUAenPhI1gUyGUIVNV3E13D+mAM9Z0WMxhpeCUFkQ3H1Rv5K
76KjG8z4UP0+RQ6yUNFKuoasohu9ZoVzK2THv1fujYi936ForrXgdB1zMHPjVafs
4Llk3QX35rFJFWZHLrbBAMAYPdP4SSRxat7oktvdm8w3m5EqYNkABt0Xa21NI//1
lS1OZju0DtxEtK+mht4BAyX6Q8MV3hamFFnYJ2hahlzofBJOKOhD6s5OieglYDv6
in+ZqkUSNqu0GaxaqkZUSAowF3045nlbmnTsEim6cBavQ1K2uIFs6rM7+FPrkQbQ
yG1xJkPPmDC2rlqZKEeQy0KJ0m40BPRQ6rSMc5f+JhOmKd7p2DDgOrUOwJuERumz
lVewiVuP3vssh4k47F1XYRNsoasS4jwXrjr+Ks+Yp2+yMRi7epT5x1/l3bbwBt6K
6n11IyOw4UxAocwb/4pR0w1J73syy0SrHAMdQwjRudPMwcQcclSmg76YiOAJJ/dL
gJJwTa2GS7vaqH4WQzCysv9Mx4CGKE35uffhRVsCZsiyTboUN0FnScDYFlpNNEXz
Am96K9WS2IrKJXfVvcylI8JhxgOjAg39YxHdFtWc/14T0UMap1UmU8HkTK9zQIyf
Gk0WrYrsFLYZiv1vLmcZvtSpQYuJeoRScP1r1lwq5pVwqDVGHjEXvoNAAvbc+rsG
0a93XLSLIwXyTzrZHdz2soh7hd4sGgk24DymzviRPLgvanqOsdnscm46brDTgDaE
ixY0rLaBYksT7BB7aaysYCo9s65UjTM+RDbE2pRukt8HHRCERsoW3mTO1mkAXxfi
O/MgjZ57J7foGTRSgKpgmhkSUxvFrYIOdVI0tUHqmCP5hS3LQCtfRaKVD0fOFdCG
T+wsiPrQsh4Qc6DyBHNMo+J5K8KwXP8XqENTsswgSTA2f7MlF+prb34GgRwAM8Nf
HlDHtSsrTkw4E5PPRvG1Msoawlz25jNhRVkBeONnsu934vme0PKfyibJe+hFlb3m
jTQJnYmCrAyUa9HDt4m1/Aq4AO9NG6oOxt1+/wC0Fb1GPhvWyiTU3ma/45PFPQC5
Zl/ICkdrwB4Tc4VtX1WW6H0kl8KZQUH6vZsRQFdEKZ932RNnPwJFC8SlO+E1bdic
5IpjwV5yC91+YkAf1dzjVdUIttoFk+wXpw0o1erh99WSINeRujh7z2KN/wk32XxJ
/fSHuHi5O0PA+JQnCAn8P50c0Rd/bSF7DHBC0PKbDyL/931J4kJm4KSCvl6MTiGD
uwAhCifywFQUhIfUMmHSuvA8KeAXyh/OzcNluZzEM0QDqZzg6/C4M9pkY96hOl9l
FODTfhns/BJ7ea18zrIVIkiAJQJps8FVQPJkXWw+E2Tzy4kCGJ/8+3VGHPcfj9cw
F6SZFsjR05vIAiyR0SgA9ERobIgwkJ0oD9sD7T1/ZynM1KBY0C1gfjiubnaA8Hdx
PJiQkXRrINYTdz8jjcE7fPlzQ4s4zaEXdhbdYhOr5LvwPE/9UF1Bl5iIEXWIMahk
uxQQ5IT9YnXSCdvrPhLRHK/KjLN+adupO1OW+J2/74qPdOqs5gnWO1N9CH+bdJFM
pb0kPLW76Xq220hYOzWyVXSdgfBuclto/VHdkfsVMphqqq1ivrEc79qc5Cowc5gy
Ms2HgGPFuA9HqZdUSzajhcU9MlIpuR6Biybf/34stxt0v68+ZTFpc8hsZDBj6QUk
rE7Ggv1XqJ4LAdaAb0DcGgO3OAc3ERe3lfaTQcMjQVtilWiXmWwhnLaoF1uG+OZZ
lNWNPysDyD9/c9/JDHht755CrNbN40cDa1fkDxYdZc2fdCP7gBdnZB3bccAgjnSk
rIsZDVG8/0tAtE3aoBTqu9iU6KSqB8DW71lfW1CMintpm9Q/5o8Kf4oyM5DbJuxI
+LsZDf938GgQDmQWBwz92trxCzDzYkPcnpTtqo+CN01QIKq6dKiIRLTFhQ6hn9SK
vGM6Im8FFD2E9ybaXvuwZ1iIcgpikDUEARN7gQ0jY2vrBu1fd5ZUHlwE1VMT6K0z
ssRc0kev7Icab0xkTkF4xTfyma4xIizIylX4AcgYmQLVC1K7LfTpI4d3qWpZYFlb
jrPcxzQwTgHiXz7f4Ln+faOh/mHTgAjMyKMloSehaONF1vgT2M7apIeF1n6szs50
ppvIdu7y2B0k5dzExyPZMnWcQP3V4/f7rGRW7f/peszlEsAS3USLpx0smKRARquj
hsYBZAKBw3nPyKUBYTgNlg474eYAEAjZr/ytG2GoAV61wpGF22H0Z/M6DPfJIgRe
b0onztZs4UCwdTIVBXM4cQOdK6xt1F3D8nuKdyRLPhteAGQy8dTqyCayoYrvOY+H
Jaz7YyCvxnIfIPUMKnRyFvaGyCFwotQgn9H7mIwwvkvvZbcbV8G4RLFffBDtp/84
cIVXBD9wqqfy1yZO6pSSSW1kcFR0IdZyK6ECMBr7SQ1X9yHGIxy1FrmjjbP9+r+k
P5ZmE6N3yICuWX4bITyZmlF1njBnktlcjlgUXLK7EGB+tKS1LE133ARpZSxsVk17
E1BfKH4bqYcgDu9qmVNR6ouBfbvGCN+Bv1CJjB9sO2ub+Z2wfaR7Nwzi54j30uiC
GY4nMO8EUYSO3TEi3HnSeujIZ0RIuUQoVTQjNmCMVqDfwHVtaynS737t+hWfdJGN
RZYIjTuIP5KA+hVStQ6wn5kEXDmTxeGa1UUhdtdf+D+/GBvE1o38vrYKXIgUFJ4T
/8vQaXmVtPXsCDQ+QsqSO0inRRno+f1hsfuJrBZYWcL/Sp6vhQwhkTom/Ulexe/o
gs23siz92Xl3V1oQKTR7Ng/mNGRQFGM+0TcoPkStjRMduAoy+CFYnjUIeWc7pF7e
qAZzfjN2oVRAqZrthmXYL+QRAN+F1PRcm3NjNTNjPbCtkQ1ouayhYjRNHbelA7ya
mhefeVct45SI+/uzKGa/Z5ItERhtF4wc1dlFqSOwDW3+oPV6c+Z/EXCA/uNppWRD
ap3QFubzFxZXoebhOEiPH2/cYsxN4nmSWLLYJDchQmqmpsVUl5Hoe3eC3ahsWdpR
a1C/x4r562kafMt2PuNX1hv7yqQvX/tskQ/Tn4NehATAwFShiYtRECVZC4+T9ZkZ
K0XcU5gBWzKf+XmWhd64D6PqKLdGWaplqoDVbNhuWYQymcNLaHHypoThRv0xfOfQ
j/okm1xdatutxGZF97YdF4yOM/twIAeIKiWwICSxgl6ZszTmaSEcZ+6Z6y5bGZSE
V2ivJPcZe9PgbApGyAkT0Ui0Qb3jtdKuPF8S9HI67h5ufmeRlPpAdkWUFGcXGuQB
nF4pMJWWHyAJ+W11XD1Mvp0pqPoyhOrsTA8DdKJQpVHfSuBNv/vMH4Vh6QtLwzdN
10hD+iIU7Yle3mzpJdw86TvmAk6DfqxWL8JtU5XbaTxqooXZloatQJKFZtPehZjC
FhUl1oiJw6OJ7lvfhJg+vNcm/wl56TQWcUacSMuAQpVN0xZPww2MUpK+BDfL0nRD
qmwMu/vDbkBdQiPz3cuWjjZiHQxeKKfzhpZOtxiaTcKYRhEaNmfZ82jsziq69py6
bOe/6YQTVcbw5a4jKKQhGXmQAnN+LgDz0hqLAOtMHi0GhwVsj4P7uL9GKOG0cuDC
LESWQQt+DFEXJHTw7dI5B6nTHwuRieTXr7B23WMBzifzAtY8n5y6fhcCL3yF8Dsp
br/I8PWpvKkpw0hyYunZ6MTaI5T5iRiV9p4OPjK+pyBn/SnOgfu8a1ab3+9SL0PE
c4Q6SJ9gKRlSAr8gXBjsvCcMVSbLTCA2gAWLBT+e/HFAqYGyXNbXlLm3Zu32jth/
dgSFr9Gtmzbf5o+6AjthTFKIe6XzRhBRY5hcBHc4PZ7L5IOlXzj65i/MEX6imEKQ
qIwmf1OUPyqwyweQQ4Cq9jHtNTgsUgoRI4aNLymVSbyYfLbebLAUOkC1eRv98PjY
7IVgF7eH3l6H39eBgLhMgFZ4M0jWctBV69ouZbZvoBxz5Vqv3Jqbb/FRkbHm48YQ
Ekfl4f1Xpn4Na3GJ5QUZ56rTuBA0hjLVVFVKDw6wuxpuSiVGfAO+Ln6k4XRI12ce
069JCYoEOuvQMYsYhL603pbJ3J3PieqTYAXWNjcRmnmpRxY4/liIHGOGfclEiFLP
DJs4fKwvyh3vRXYz7j+aZZqhzM5379FZCfFVUcFtgGgt24Hn1EXpZzH0i4X0pKVT
/0Ah892ZhxZBTzbXvH7Ae4sIrI2IzNVutj4adopjSSvGrBtoiJ38mFTjpHLzhc2b
pViTrzHNa6zKCMmaP59YpWf/9k7BXTohsKq9CP78XC7oTUV6pfGFDGRxceN8cIBz
4DtQKa9PXFpLP8PF1L6MsuUPt1gKRxBZFPuCKu6f7wRMXG6AHzWBdc9xaTH6QOop
i0jnSIEc1hmqDBIrPvm9tO2kj2GF6ouMWAVxzgjELznZLhofXRNj7O7lrLnTpt3i
DECIBD04c5GtYaMG3SPOO4oK295lCdy2yjW7pfe81Fw6DSsM8I3JCZNuzIqWompz
PhtknR7cAcxG8TnFxjSEYK2OKDnezlKDjJzx+EZ2WDlmW7YpJj7+xV/hbvj2DuTN
SyqV2WwWeP+1LYFp/DF01hZn9P/Xzo0ErAS0xIElR7/fAkT1Niev/NxCsXXGcv6/
sclSZTDjZxVP0c6w561+eYBIEHDHjHNyc0QJ3BqfTYLwRkejT7v34IaIjbEkYvsn
JWSNz9IZ8wiy9isOPvVuPsGUqr6J/UJUUC8BrtjqMP3L/RoXk9krdbVUdrHBhcyz
rFlYBjM0+K+eAeXRXT9o+GoeSUqW4Qp1StR3/oDZqzVV4lhA6dOiuGVzHmNG49+C
U+xV0kYDP1HOxBhih09SZkqatkSUHCPdfeP+ifGq1h9FlFwPlDhYi2Rx1a8evV/j
PeWjO4Q1jxfsX4LspIgKxVKN9Kuq2d3S1SDLO4tBnV7JLy6CAgTX2dsXRwu8CGVA
0R8ff1SetbKuYYDqJ0GMYKav4RmrHiUsdnUhsw/DCk9zVDKN2u1HtLtUYkHcULmx
rMpCe3JFuSRvKpLwDXoh18dJJIKC2vnL7Z4n3HJboCHiIV7eo8wM2mzOPmxAEkcG
OzDoFulAqZP75yGDLwXbygjFBcn2mDhD0EWcXlWS+hDLGwXH5j2cz7Blyjcd00tX
AUQBYJET5aIJanXj3RsZQyvWq8F96fefuAxzGMzh3oUOT4UpywdmeYYoBi2z3Ak7
evPTyOFQ2wrI3kQvzL9Qz4trH1rl1krcJbdVS+EDlCOps7m38ve36vtYJqfF0RWK
jixAueal0QS7//dn6EylxwsEk3qi73EpIpwLzowMhslzo2LMXG/hxxz84Gw7s1qv
JzwJcPLvppp+lDMhFJkT6GoLasgnjHyUZRvMG714kdqS4KmUs8CpGtiGsjbLlTRn
QakYa+oiKdJykD45PuzCWI71I29trfzyWYmr/+ePQ6rEX75vdyfc5U1cQMwVtX37
gk5xQ0Orwb8CaBOstuABavXtpHnpBZJlFbhh04RJvJj9u+13fwG9nJ8FR2/WTqbV
64ntAihmSOjWH3szAwsfZH2ngR9SCSNSNBJFyXyhwGjIXo8Id9Xg6eu5h2mP+b2b
idFNqDJ/UPeFvGXfoBgx89jtPn6oK6IL4zokFCZv69Id6W6fBhH7752xdm2222NE
t18bj8qHiue2b9yBsBcbdrVLCh4pcj/sLFYJm2JjdSJb+Mr+pOQJ6KFQVJBoT1n3
kFSjXnTJWJ1j8HIzwT1e/dMnV2csyAPvKMf7dGXlwDOvd6UqLLl5Iu4nXXmSqXCP
v6yDkomM7zI8k4tYfuZzF0OSG/6tOmr4yzGxw/hPr3UFqrEjdoDIki8zFQBDz9J6
xg1HvhWDJlqKB1FhtYUGzClNzde2fcqWkQ5RDd71NmYuLrVrorfiZJDl6CDaaxbA
of7WohyYUCkaVfD6pgPMA2CumklG/O+1nw2T8HXabMV6VPDkIFnE4q/qZVw4HGo4
AeH1A1BA0uH7LGbzkFexOvwkxcZJbGVW9D4fXi5HE6E0tqseASKsfhplntf/zLip
ZUCkaDJDkdOn5OKj0pwO/JiJlVKWb6JSwy5hA1BewcuHaTzwy3RtSD/UEwFVKkf9
3dm7S7n1PTIlLUPRmlOu1Wv6sF5c9aXlwibnSxm1X9azAeOOFAQHeQV4rvgqAlZW
sj8xkUym+kySpBwUOtMEEwQynGyhJE7zcD7ISgYYfnTe+vyty+1l2lfNAQz4ttLj
9O7hs6Ri0wNCIUWhMgDRaHtC0qwN0bC47+3srbEyq8/z9HxQG9lnLQjUHBBY5CMl
gFnuzW5bMqNvOeu7jatjNGkTXFBKLasJ3Uuu4GTk/x2l9aXbRSDNMPaj9WsRM1dG
3qACKsZRKcZmN+8aI2pTK8kPy/D3w4wOCbmgOzymK+qWGBOYiADo88d6/xZ6wTsK
hBl6haZBrn1UtKVKEOpLPugbAZbtNdDZ+Yrmyt/ji3oD21acOGExuMShDRUdFZGX
yVeWFeXrtiCBUQNe3zeQP0cYOnTxVIWELTTZKVZeMtPOZV88M6ljYI6nahpJQSu0
I+TQpOYEH4TOcssbDmAGlwnKkHSbEnO9Bwx2yvjPkeXz6fomvlu41qrm4Ca2HgXn
dLgxXfyeHoVLlrEwMVG9PIHrAQb9KN2kppsx3xSnlf7YF2QLE8qjQ209RwTOZc14
neu/XvDLagrnDWavlqV9JClbYMnWpziPp+uSdy/9An2KN3yLv7M74wM26ayCKKWE
n9i5LZE88GuGD7CLQzoAEik7OSp2SyX3bB8shb6a6bDYoUfAPU3tJX1OjBfficce
ITweIo4HJRKGvCU6cjtRUUvefMevgg6DaTB6lYqrZ/kPPSRORPslLwhi8I+P7uiT
wWvC6ijG5kombTqnsGzthGLYvZ1cR0MfXuXbgj5uharZ40Nost+UE810maFXxTZH
IDqreZ6a3zZg7eQg6IqCqqHyejYXe3F/7JTMOLekzahyv8mWSFeXnd8twbgiqB+3
qO6qppOomnms8A0nUxg/lI2szYzrgFWiK2CyY/P2jwJDyKwGkLTcsGqVygsTf98p
kk9jVeTsDmo9tOzq+ABr18OtYqdw9f0BBlIJ38hJ+HU/ArlFtrnwFhr6qWw/eu4D
DJr00ikxsIy+CoERIITizscyNlRGkvHDh2CEs3zWNlV3a0VgLUoJ/p+D6ev7kzfE
Hy9Azb7MHipAYr9RdhRQphGEtD5OVouZm+Ym/HYa1p4RyRzCzEfy11THpE6CSNbH
Y7QUYFDmEtuToq5iPwDhbY6eid+nz8wpQmvtp6waVydotQmkdKFW4Z6G27Tx8y/N
d4hX27Ax9iRZyBgJFRgg97D/qU4lme3SzOqmbWW5VBjLoxszMI47oH9TNtk/uINT
n8bOvObE246GZwII0TbsKb12RLmOf/TrIxtVLfbkuyyQuRzgV6gcy6NXLdLBcVyL
puQzNvNru7HWH0hr0hyM9xfio8Wek9pqnOfR/j36hLmk3iEiMuuGM9Z52oQ84sl8
rsBWxIY4X6wy5FaaQib+fgH5olDVeo9dY0VZ4MAG2aZYvRMVdbQpGxCtRwU3+JXH
bF+u9Yl+v7rbBVA2jHFLYAAcvpQh/boh64B0vS6MCrO5aDb750kj49Nybx1oithN
iXj08BaH6z8p49qBnhNEhgCChTDqvrxd8xf7OL2I7bAv70PMbcPfyR7SU8W5O/Di
lok/KjNibOzBDjBR8qPFoOj4SDiFEdUNre6zQlCUMiq0jVaD3VOr+wIMrN/Z79xE
nZVL3EiEmvMTqkaYlhi2z4E1vCRC7hr6CpyBmfE0LgSlEd2Gt8m3vPKoL1nfknxk
wha6vSPT0EGXz6y7Al/FvcFOjQY2dhC71KGw4WkZmyxOZQyU5xt39lmQLvfWmF8J
qztmEfKSBsjsViNcRmy6aCimOLCnegqEeHglq3uvkYBENALCR54z7iZkLDDHFgb7
fShVYXEQb3jw7tIgAPElz9Inpbz+t1Kvfst37yPS+KLgOkSiIMqK/rUQ+yICBVPA
M7PnRbPZkOdZ+tBA5E/hiy3/JGzYjPCXnBbO7MhQ8gE5gwKAPf6EKJPaHcNI5Kk6
LQOZSVZUUsvNx2d7M9xRbeaQ90ZQkMWhDcWX1EQUdPvD4qOWX2U2UYhwCAIjDTjq
DbO3DIWsbwP3CXJAj37/eZY3yQ4xY6oEchZe+ugeshQrAnzPuOFfkg7cjCl5Wg+N
13XOmx2UjX4cG1zK48FliJmFlg4kuKqzuCsixjPsI4rwK5DsxL8JdV2RiZYPD5dK
D1YYx1MTwEhdITfY1BOk9mdOzS0+YLlkBj0nXE7g/rMaxk4Kwna5HmhshlWtPdkB
3yEIveQVvSg19l4IPInyewlFsZ4Tyo8ra+j2eF8cTerbBnmbOMzxmTNPkLaU9D7m
PZ/tre9CsoVNCjtbMVi3wDWq/CCrKYeTlJzYRFFtLT4UVnAwtrJpjJqHXwcZHHBT
DdqKD0dJkbxjck75a7RmNYhUc7AEXvsT+iycwBowI+5uc6s9KTYo7JQ4OB3NGQbp
5rbl22ZvqRzzOv4Ihbnkm1yYzrFS1TfiEfyTbr4uYp3oIq8JsuBAYbIbtoyXxlDS
4mW4noLEDdCQOTAfMs1S6O3oLHqpY0nZqgr+JlVM0zL9TSNaJ0d+ZDrgh8MjHiJ9
leY3ZNth0+SGrc3B3G6hL4PERarzo4T0NGcct4Ex0D3rW9EDoe9yB/bhejdHPpEr
6ZCzFxgNoiMy4J1iPH0AUZy/GKUQdKP971VihBqz0ajZ/dUYnJkilo7qQuEFXkAP
4RdaQS9dFthL5+jXryZsqplvCrZbcNqLATh/j0RK43Owu84WR2l4l0I/aPPW526U
HeJFWqnawvI5zNA4ZtLTwbsp+8qeJuSONi3KrUnsbVZ57ahozNVtW0zDhzbz2TWq
uI6gHe2J5k6njajL+Ls/1SNGPNkN6cNW9S4pMFAM4fBVPNzbn+lMDsIjr/mM61x4
qrTlPSuan+m46kC/1/CeqCStWhXB673lZlC4brXwVDaUiOwCP92+R3pbR371CSoR
o276ZEmIgeo4Qo8JFyOmY8j4+dw5Fhh2ARmxp3gvdipC7P0MMyc4lECxPss8nyVh
HhENZ0TimAD++uysTVqBru9UK7Ku97b6N2IvrHhv2z4+336Hr0tT4WejrVRR0e98
xIN/4isgkY7FTVsLHM6Klbw4Mx4yh2Wo7Vx1Q0/0vz9nHz2HnPnqs/mw1e5JzvUM
eF+XTCqnTcL9wTEhSJtCoY8mqSSb6B6do6SswdrrONJtOVIc5NDNSxUZ18t0dAWW
y/m001KePvp++IT+jmM4aopksRNBhvjdQ4KzG/I9fNn4Fp6PRpTpJvN8SlgDVBxj
S1H+RK0B85gAXzh40ErDMObZBu018SEjSvvTQ0IIQP8D4UCKKvr2pdgItLoxzLFg
ox5OhtqcsaSDmrvCv/ptnfXqkp/Z7NMz0QPfLNk4WV7ttk8giH0jnVnww6sqZB1C
qyqLIhiMHHf9mSRQb33ZL53YbxIc0A1jCAVcPfha4+rRVovYy7FK+3Xq01sROXqU
arTOYoEEX9Xz1Dt3rWyM5FCBoh2qRqIOhVXzUgA6HlH9KJXdrk2j82EoRn+Qq4O8
TUX6cD7QcKcwQ9wxC+0Y1UUIlKcV2Gls0d+oFIQaqEJWX3+709bx4bMz5tDf8osf
U156dXWq2mLTtALth9iIhXN69gJjrV7LBz3wX3xYt5TEQe7SMn0F9rJXlRfweGZs
l10LJ51h4XIlIjYq450NkSljEaZZ6lPjJ7gBhIRAny9o3Thc2mCyPjbD5uGYBbl4
6GJNsVEvAYAqOGzue9Twncra3XdT2mVYGil1CTV59WCwZA83dureqpn5/GfPTKDC
Q4Fwi+EitUADb2H/3Iw88aBhMFATFPv0LYgs2Wt3rRRedrLjBvDExXgQqF6X+uqi
klBuLYuR9M7JRS0RsnXtRXgcItMsCJciHkqXWBG4CrHTQib7qKsV6MVlttHdtCvB
Nvn0dGUO+VxXmop3tIPTai1dcMpu+9nt1P+LiVEZtW9rgsxJzSI+MQ1jUkvaC2JT
luij2hWCF42FD3mxAQroKEkxS7Kr/pq6fSOA4uOKswGkhUWrY8c6Y2W/JpL0YqNf
SXG1uQqA5lkTWCVJGjHMrXUce5xFcTX8e4yCqnUP1vM2yDgTk20qvPcf0Lboybee
wmdR7rd9Z1JPkHc8FKYqA8rmRFzm0HHHxBeqF8mF8ovGudJIdeH2bvndyH8LR7Kk
sZP+4RTMk1IvU3o5SyevfzAsVfzynTVkZS1kHJKCLd2S604XR40RKwdFCBA2yrt1
wfeuGmSpcTyVWorvB48hQzXjMda/d170x1L/UfgntLjeJxUkj5ncnFko5G2n6U19
BFoi0cfIymsinW4qB/1wNyBV/hKXURKm29+ialmXbuYUhYVPMIXauxOs+lAq5Fy0
cs+L0M9zRLS7HiUq4PcoEc8Uenb/JIfkIa+Do2MEl7XIZH8C+Mo/ympC5Cixhjlq
F3WOPz269HmxVTEpfgdfBtTPL80Ry03Ev5RewXgVT9qAzzPNWSC/GFZZ0L9uzkbn
hcSA08Quv5KB1RCLI3p0dPm3h1YSmpB/d2VxAzKJZuMJCYpihE63nxOlL9Oytaim
ORBuUQOZYfgd6c0nr4MLadbDO8+8M7eLU0JJLZxa6vk26A8aBmyxMSfTpeSNHXyt
RxcbRF/fSzpkm02StR2vEeH5vZiwsjgCq2PHgqlhj4L2UT9vWOW/BN8NmVOPEXdm
Ngeri8S0vMh/iWPBoEUiJ0Dw+aKbryMGYaDV5j3f34HUiQb8SKwm2ZZby6pUA2ms
Dr+w+S6c3D5a4UbHAPQA3/eXE/fR0TUBCGiBJZ88ssBVss5QojhjDnUhqmQYNCXi
h9NErPqdH6g5lNh+DMuKTyyGO+pfbFZ/SJTLT8eHEggocIb8jq2uQY6OSEv1jKA3
33gaQoR1GIzMNkgaIojPkCB5ILe3lkmJncMkXNheahsrEdE/1NKLF46/l671ifUI
aCpK0L0+uVhhqRDErZPb38sOzuC1pXkFJmuo3WQsW/AZ/+PeAAED3Ce24Y4fGeaS
U2LaKeRYQpyyNj9e8D/ieeURzxr7dPnSjS5KNfpbARVIC9CJS2pw1h1XrMUVOu2O
LIvC7vU9bDZLvo5DXFHAGrurA5OK7oo+RuGhzkh1wbcufybrJ0UCapy52+UUMuCs
CY8kmL9HsptMk8SEu0bCTn6l9gx2hEes+nTTuu2/Q5TnjFivd/eA6+vfT7tEpYd9
2moPh0UZpc80sBj8ACjNn9vJtW6EMoTQHngydwHN9i9FD3llWwFV6nLAmc8UVYLE
0BC9+6A/1p3s2CL7WuzovlnqmvdPUYOrh0yZB6qicDsqA/B/Y4wOW+NGBmekYVpZ
WuZIDBOl/DZe85ATHw04YGHqJwh0CYx3zPv/SSxJb/ggU5vLNUl0AzhpDv2O9SRb
Bx3RR2VOev3gG6iCppVe1EDUzXtJjYpSpU8ejxFQDqQjRgpgEZAXmOXYv9bg14Sq
4P6X1glJnL8nm5EncN9scMuUgrsAe4I81hqaTfG+EL9QeaXaq+XUg0qVDuWP2wYE
mDcnqdmUWkYOkCfN+4fManvdMfJjcYQK5CJJZpBD9cfFvgNauj6bUhHZ6nP4PFca
5nyFL+1Naxb3G3IKeJnFSQyXuxkYqDlqVdi56ci3yVP15ISlakW9wUlII4P0Sq7i
uUDp7TN+7RrsPKUPQvEntOduNJnm1BytrO3VaErJAo9TYHH/Yt351Q2JdPOpzG2V
YiXcWrCbdp3uuD3FR3rwzt4mbVmyB1bUNcNHYy89fNltT0TIpJmWACJg4Oa7+C2X
RVKCnOdD7ShE/T1UJvqWMU5rLs65pQtv9a1Yiwm5EW+fVTPSETYcR+rixY+l0ZaM
E72TE5b0MtNP8pX/wVVLyqdpjW5D07WEfb2qAbmZApM/TN34uOx8gmBJSDxGWpBB
R7hDpjFzGisMsBi/Co7bTnSnQM4RGDWnhTswZu/0188tBXA28RYjoV33FsdE2y8T
a0v3kYgNrhVlsOflPrHOGbJk/mX4IgUtQLfDdMr4X68wN3cIS5ctfsR/HStBolKi
1WR4V9z7THnMk3d3l2xrxjuHPNxaUdqDqEeE67VHC4XWoHjZeQQBtx+7H33yf/24
KxdldSg6i8pCYw9U20jRujQOChpXRcsyWuxAKPhwcbwwJziLC/kHcnHRtDftKoDZ
/Ib4OrHxbXam25kjKnNd4HUb8tTSHCqBjdADjx8pqXly5b3HRo0XQnVQRPUYFXK7
59z0fpirmcmSLbQDyeJn8SY5r2NuIAM/NhikD/QP1VOE8aBz4CSo/fGE67184W5F
gcC9bJ2FA1322mGAim7Mvb3jvcmM8LwdPGBz4V7Bbmb9i/q/bNcyJxdS9GychqX1
DrrYdh1AvjzhzjkZBZlpPPI0ELU/QIFm9gMBUl13SRz0c/1tZ4R5RLt6liEvZVt7
egpDfQK2Y90maRPOellWB4UeqBvAb3NjRgvN6RZRLCiwa8G7X9FwMbGicH1ZTJAH
zqcapV5fe4VG6FiJpnDaUXJ7gyuGObok4P1JYO6o4v6mFYMu4wUTTYS/HaHConoM
bTt60Uj7bg6lpvXfvYQVeblHwHUd8gs+RIFx2wIwtQjuROZ6k2pAamSdJXCeSZlD
MujUEPRtl8fViwcqbeYfZwxwNSJhdPBH+DJ0uly6oKnNYXvp+g7f/8G94gYuPvdw
6r2w9WP5WsYvxbqJMIkbWHRzX8Vdp5jQhntbMd7ylpN12gnwVg7WnGpH9Z9iqSnL
GfJSpdW1fN369JG9BbyGC2P9d/9Gm6+DDKvg7nLsbHZokFM4z98K+mMStj/510xQ
T6b/wDZr+v4WiSNAMfwtUU0ca+tbvt0ejDGt3oQQx4Jc/zxyslBPzNCIydlPUiUW
sS/DTtMFI//sHMTc5PQzCGPjPDkxmudIoeW9pBWyp/vV7ozH3OXM0m+q9b4I/PZ4
YSa+gICW2QEJL464r0vOi71PJ36OrK21HDsX0mOVEkusUq6fiJdILUWV9c0bhIOV
liFqFVy+mcldkAzBabyODI+QfbTgeeBrB7fttE+aDSroEI2AllZwjLkqb6Gvz/6P
6O2LPeom6ioGQqpm70T7dickWKS7eodKUQK8D2QCngM7N24BWod8Dbl5swltfyY6
osXS1jcS7DtnkO2dwSSgbNqTtkaDSw1R6qInPj6gXTl0eVzEfWlL/ARzIKDEeVuP
uMEF6qmtu8UEUyOnlCj/LhzrRBYqPCrjOpVnZCYTDbF4LpNsJsy9ZZmXfqOjhek3
YN7FEfl3HJ9/5NAgfmadz8E393b5VJ4WWdV6VKjjEKdSpLSB/lUoWVYsJ9Vc480H
1iaxgn6b6TOh712XQzLmsjuSJyYvCSRTqO4maIVNBJn4zBqkbjX2L9AOCrLyJ+ou
ZayRNkCBh2aREjI4LhlesWBqoS81CLwGlqFy1PpyK5sjZU0g6yW+KqWy9k7x3aY9
QYKgZ2imHS5s2cqdf7Twp+KlQEI7xSE4nT/i8khgYidM0N0rKfklmOAlbwOdEHA7
t0WiVmUMuTgfgUqvuxrJX3rm+5CCNj/PyiulSoiPRK7pUlNlKoEo7pt/yPR9nUL8
PbHcXsGq3F0o5+AbaOEiTF7c/4WbyPwz+P3F7QOqkqTokJAIpWHfUIqwGdq09gFp
RMUtTUMkB3W4a1JD8GDHM4phQftkXgUgv9W/Zg8rxbXRc2/ik8wBnZFPK8bD4MKa
kejG4ww2cKdcR/nlPtzRya47kTrvem25dOE9aoMmom16IIwbvSBtkH3aOPHCw/YF
ZYOAqNCkC52OWDsSGI06jajPdlm+lMTN6ZtE5qlzDNyObtXzqnU9HmqQPK3Ri4DX
AuwG2Rc09cVMHBmCfJNlr6Bkx+lQu/c04/9BEFLO8RDcnihG+UR5nAi+AIHpSFV1
fkwSzUM/nlj6NMddapJxf2k/fyEUYVgloW45o++TXstEKalDxQMPdtsXq7/7cHSN
9QJANISQrSC97R39FcQ6t9k5T0j/glT44cT+jcTSRZmbgZ+PII2cOV9BhJNndrO/
/Gbwk4KS0wN9aPDoJUMSfwDhX3aTzPqOZCmgLbcRgNg0KHs1+GCM/EZdFCOkPda7
CVgrOyhbQpcYgO6ce4zTg94xIKl7kClTvOaUmFCbK2kVPbHAq7rGUiXY6qvU58UT
b1nmWjLbvpiEfalSsLhDacNzpX04Nsx4Yo0QM8YZay/gw0CUJpvK/gpcvvLkOuiZ
IxVgIT7IV4Vo/A+935GjXnh2fJwt+W1UXbnEXFuPAGn1NqxNLLGVzKxgyS0+1Ugx
o4sUxFnjEUkEuzy9q4V/ukxpQ3rKbWWyMn40J/iSWEuxQJo71aqpVMGJCwil1OhM
A4ywGN/YRKg68Jfq1Czsp10i7VpwBpDWt5V/ZgXjeamqxAQLzEhGFrcLoGjD0gsN
1qs0qSNnZLo28R6Gi1Vwbwc9ROnIVlCIrSsDBd8YiYoCZCg7lkTRKZbMtjqUKkKR
i0UY0U6xVJ2BEPVUnqhXpICcxX1/vfeT4d+Ugi7m4zRWRHlun2k7MMQRq8ngjFs9
pS9aVFRrfjMuBTDt7pveSPDYRCPL8ndh8KWDjk613Kw8FFdtxIZgz+NYOl90ZL3m
4mvxtfVnI/njssd9fRuQThWcKiLXp7nh3DXSQfDNl6IePWoPQJfeXNWlDS7n8Fks
ngFm9zpLK+lva48fIwJ4rVPrHqg07wvSRsyEsmj9FMPHlnhPS/jnbis3HVft3Pvi
+7+mDsYLWj4cZr2/KrWWXdEmcbLhssRLsXOkFFPf3nsjGrscgYlqyy/v2CaGe4s4
Ypj94qIpwQcAwQmuSLHI8Xm6755xJIWGizNApR0n6du5XbHXlk8RiLIfUxW2YAIu
SGAsPbDtYbdaM39vEbfyKgKmblv9IaVBkvpHoIa8HPkHlac7IsDRULECGBsCzGXd
XUsBrHgOoq3da7eyA9sQ1l1/V//t7ogFhtQr7VbkRQ/ujKS/JydTSM5lyEnhuT1z
RwPP1OU5Ipelo5kb+7E1q37GBncuJZ0/i8rsrXKE0If6rhuoOumf721t6TxuO5Lj
o08e4mk1qB92f3BZ9F7/mpzjAxQhzAKQcvJYLbemyY/I4R5250iptHx+yOLBhiPI
stject32sisLQCIq0+VooEIJkhdAV+C38qUEBBbWhWNMc8wkjkvqHzYh8iN7lN/x
MDmAd+QAMZtJw0Q4+yG2A3eFeQMiUtcJrkK1K1mTx8+TX2TvTxQoiqYxpy4jcUx8
vyqzJxRVjC3JoBJIpzhSz2vvbw5ddICYrPK6r88I6tHANiz+QMatgC3GTQuQlF3F
4FCUq6Z2DQKllpD40p0T1wSxnC3c/MBdE/T5dTgAxYXqGoQycTYiwCbGwELHWnJ7
hInlrJYgBsYbSTz17APCupNEBIuT2t+pFDZ5MJcATtVykHp2vlkk4WzuQ5LorfJa
0nNwWNzBjJOw5YV9AdSlGSFeY5nFFYtyMPn40hU2AypkTHVwwcptxDUOCIkhIt7m
c90VJgtuS87lB23riHmUzBT5+khs0qjliD6aFr3HT0EcYatXAvmAAeK3jNZl1q+X
JNx1yPOdNgxHQw8h9BAejpbjuIeWWckVglaijSyEvtysP3vmR4JN/QkJjFdCFupL
3pt+nIO80UuU9yeKkiCYm7DhDhUkLoNkEVLE+S/93njxr4CT3y/GPtDk59FuTwtk
7WyJOBzNUykQL4PuXLsTilBhEA8DvjQxuT8B69tHksXlThiCv3REF6+vhdjVcwlV
1u8FAxnp3f4ixzCrtvQzYlbLy6FbTtZUUPozpz3GMDvAbgm/owmIHVEd+8Tdzxoa
ap+viZEl0jwGLl4t6LdCCXqsqB4uDZYhKbEfCKA5HVo7OEcKGwuq3B2QZj+0xSVv
zRsPkpEoAn+Vh/Ibjb6gSdRBQRFxugctGczH+wS67srGE3lVXpF4tiajzcwqe+ih
+yq0uV7WSg4gw5SyDfDeXk52KLCKLfhGjzfNTba6QV/JC+eMYIcRTJpyVycywKHG
BGULHLhstFrhepTdVl8P4uHYJO0PYICYXAEs99MpRDemJla1XFvuoHBrn8qlEOL+
2Kzdj1LFuCIFQ+p0EEoMG/ndQDKmzg/jDEAX4copugHeIEEDfnmHjdE5jr0GHEG2
nxNbIHhaHPFSmbg2/RjjpzqNCluBj10IxjMvgSPF8g+KLW+9NzoRKiO+XCnq4jdA
BEmxdiXCkgYF7wmL4nxqucJ4ocGHCLVJNCmpM7KF+kWu7FMe9W7u5Ithh78DDHYS
7dhbmgo+0ug2gjcXlkyOvPpbTOJAtVtZUdNU8B0x5dKzZfYGrHOGBSq5g5+z3zVG
zw/Z2DXC0o6IbwVbKmSe0t2nB4yLAAUee/zzAN1+XECmxW5Cw0ovFYwmaH8qmf9P
aZXrUyt8CG2Rr8WtxL+EIhQ7i8VzD0KbdbR51KOiYNA1wi00wCevfDtagAfJGZd3
Wr8DYhQ3+KaqUC7x2j2MRhcMe1SXHkuJkAwyKV3ER+YZ1deSFhsNkmeO1l4K/0RH
PvIItgckm2Uho9j2f8a8B6F76D++kjyJJY6SKwWlvnN915enCHLIdD5gO1IN+Ll9
AGksj9aHL3NRj/0Mr8dSNgkwmhY01l2Tj8mR0svyeBeUtho2sAYrKLG0FVZ8Gye9
dVPlxN+QninbZC2Xzrq6aDlGNyQOKNLFFriVxXuj76KmAcTp6ZrsP4EbZtxFSqoa
M+ilqOLgBNjECYc5buFjiAyy4BQms57wkfARN8FthkcpBBknkJu+4xxt+Mku9Shl
ECbemE6KwY+pziRHCWKvvYUy8ULIBe4YS4zWIhTYIv2yfVsS3FgmZFBO39kr51Xq
+5fUc71oBca/7OUrg147UADHGMp9pK2VbhwD6J0qzgrCwr8P3NGM07+K9MiAdK3C
0mpAiwCPv9pqh3hfwKrivwcuWWAxDdR1vG7nT/SqbvAC7DuBlvxZgYRsWUctuJB8
TxPk9t1vrcGg+UX9WGr9IjE6L53K8fLzNC9YAhZzlUzPan9iQFOEy6w2kaQKU9Lf
UtXbelZbOqYBeIO4TLzgnCY5KiIVz8dcTPPCBYs4V2XAzpedPCO22o4iTmFYMJbp
xpTWSSb37mQ7qPGkZbf7lbkmIfX6o+TOP3zBF3uhR9Hp9eGWM5QqSdbGZEA91Cuf
XQLBztT2Jj99mJlw8dtcX1VwNIAeDYeKe/2M7cI6kznZ9pl0ixiiKejUhGr6Ju6O
R1LtJHmE23JOWGm5+RSQB7kb+sCFsE2f2i/UUGRsNtE1lkT6OSwC8+ZLvw5Atn5K
yqmj37jp0i99209XS83wS9uBYUFvFAOlSg/m/fcBGnMvoXg8SOjSgAdkr9AO0PLZ
DO9dfhwSoKLzoVYtSlE6vJuakTCB+EJT1bN84NL+hrCY0ND7fsilGMbhugSuP+2b
HSiYLBEMWDqeOHhNKA2BPzyP0nlONm3Gg9oOfk4K+Nm0MqqRFJ7c7HuaAflY+rv8
zzdm7BFXdpW2NrkGvUyNAVUTEoAqX9Dyq/WLpcY+xEOnf3OwPaqE/RogZz/gSmbx
rHTzlRacyyrS2mpojQfA2EDgQEKfZUCE+1fVJCi9tNUGixVPYGTEcjWJngpgf3AX
HmVjuRD9StfQqeE8fl7mHJmv4Sjn22LamUBNVxdgH37XcMyydqgurpvw3w9wy+Hv
otp1vIzOa1J53ZOAJA6XWzu6px/JyO+Kd2pQyb1VPX/++NqYsDypWjwD3bi92l5g
VRuwgWqkqakpVJ8XLJnc36XzA4WOs3gFrr158hpIJwXQ2Ntg+5DNJwR8oXsGRkbJ
eJEwu5IvpqVPlBtpnlkVWoz3RmQUimuqa0sRm9LZ8wexeOQ+1mcXgj5S14O0mTLh
eFYSvgZYVnSgKpvY/oLrY43K7L+vyC0fZ6fuKDzOBnIfKYO1fsCg7mv+nwI9QSuA
Z4qeGmla3AG4KYEZgv5LyGppUACjz/nQPNf1sQIz5yKjsqCyEPLyndrwuJ1/Ctsi
s7coJcF1p8rlUQT1oMswBRQtn8FqugqW5x1WzQ0i7vWhq1hBA3ak6dItggD99crC
YedMO4xN1VuLsGRIesMNjQtvGDvJ2W3DwUDn6HHF9hMQji0PzfoJnf01VqYsa5mW
zNdOO/4Po4nvbYnJhZwTjHg6a9KcS6WD3IWnyXO+SUPUjcMk5BC4EfcJFKTqMJgf
IyQcTcUisSmDeBnawq7scE5YPP1b8S6YXmSadzqOlx/E92/HBv60LiHuDyXoAaBF
mVz+cHp2Sl7t5ePmwo2JiSFYdIg0o1ap7j3Y1XR8R2fNjJTb84pUaRwetZ7l/K70
3QGST764rFF27tdQBBDyoV0HuWg6XJogIwztOn7B8Cg1rAGrNBeGF2GV8EA1zRkh
kPOm5i1HAyT2B122UtdmwczxXnPHxngbC3qJYrIq1CC2FQ65PftGzFtj3qwm7n4p
NzhObRNvsGcOdEApXNDQQ8V2k6RERA6cY9fi/7mfnMNSK6Lw5FhJuHdj/QQrZmHa
OqlAAMoi3l2lhG276kd1hVu7NFFgzJiJzhhwLxoKrVTT7kWC8vRzZzpowpfREYSm
xmVPHd3xvsGbx/ZYRbb92NmUt15qL9t7Lnj0WZhTyzQCjexA/m08z9rYqWKaYzpK
WUrdat1xWJoZuN/bnMMKRXxWFj3119VOnTZ7IoGGuP9Io0vj0XL4E2y2vhi3eTIi
XdLZjncprrabg4L6FaNorg+o7ly58yrXLNZvIqJ+ZLpyk7iYjjkPFX7X7A1sS3h8
rkHmod/hpGkz83D0PzcJY/LlvRx5hNcH0GA4Yn4yrKqmJ6pmZ4fABLo42B/Y4P3I
zTPp1V4BNeBdVdIXsHuT4lNpR0G8eMypx88kfgS4eg+6hqNBy80quohRwIH9QwRs
SU+LH9W7ia/zeWQ/fjXk4Jifxh61qRiO0WD9EZhSU7EjXnaI8iK0C90RmafNcbS0
iAeGMQM4xrz7NsquDwWUDm53sd8AdoTdvwBqAqh5umkiKqweOVZOCqmskZtl0lHw
RS1Dw6hdmwpkGgFyzN/nl0ZKowL5MmDSsdyWk/QCVTHu1ku/n5bdN+Aipv9T9RcA
hZnFxwZ/3ItZ08+v6uRAmcITZoevLlsFwtU+vEsvM1xVe5UmKmazupkvz6K2yvR8
zq1axtEnKmj9cufPNF+Q7O3RIh2JUSw02ZLVCmJ4Xtva2m8cajlSptwM5H2bhHVp
xNIMrx4Fv9cqIjhSr3sGwb6zUgWjFW/QDONsBvi60sGseb7MX3CvzDdzA7L7xVe7
W0MJbOj3NudKJoPVp+YmHIsplP/HiWfbIe0Hq0dvOi9pKixW/Z6cHozN7wEcDa6Z
7enKsIeW+Sb0AwxmokDmzuwNaDPIZzvHQl9DDy0Jl42F13AwDhd/beBusiNX3QtD
WvgI9wXOfkGorSXlIdQLBPpP7O++34ZXjTeUUKaPm5qLzOX3HjgaBAUe0JcmTqa8
PAKhS0v8P4QonQm2LYEQE57a1/QO5F+lDwabCdkHhQkvwL6vvLp7HWkkWqnnYyBC
d5hmCicqntsiwHKCisBDp3cu47uZxu1jVvUoljwWbM7qAPfJU7C75OzPDetuYfQL
IpleiKDkdTNxFYlSvdHC/Zg+AJM7bXi1jAWS5rUHJ8LnYSyCcT8dhA8+oV7Bukyx
zfpFwARlLblg8oDkmN765ilhCcXgqr3nSMZBiJSXHTITJCBT3Apb1Iq6OX/FDTS4
SHHnfBkNjp0neFg5HTc0jWCERBvE8e25gUACFhNtMvP+yeAmR29gI/vJrErFotpa
cNV+m3VtO5G1iOJRb+KLHUWIe63wyAeDmLbbtNr+EuEkqXwf3SYo1x9IBsWys2Zv
lgwVflh1t40oBQtHMnCBzv/g3t94i/ZtU9GEMe/rJ6av/oqiKS5ESwFdQ46gFs9n
uXIvuWpjVaALGTPHM0ztowJxx+3bRpbwI2tQKvdKK16XOVjQegEU6EaAVxnAs1nh
VrjJlOH0FUgW5t60FLbba/ujmh8YJcNKsm+0libEl7ZrSII8xOUSUkMMK6cibCj1
6CrFgtPg1qPd5YH0Y4ryR6WL0qrrARujNNJM5C0Ddb2EbOSU1ZmXorgFlDlglkKZ
ttJLcdqsjU1+VGsT0esWTh2CqVIPbr4BKvwpREpq5BO1BmNV5q+HidJG7w/P5a1+
iJZYmZqTpDkm8UD7+bKHIQOJG1x5w/ZOXv06EmggmQmm/BKxQQ03E4RkABqP36Hn
CStkjuFQUd4mul7M4O/l6ecqsijRGBW5/THaMP4lkImjJE/tci+hHu6jNAzofcCZ
sY4IyTfPt3+L7cS+4graHlkFyoJwgwGVdQySmJnSXKYg0gUgV4soEgXVNldm/P3b
q7J4EF2h8WhpB1MkeyVWBdzqbp++fUYUtDwQxp4tw0l/VYvi6XyU2PAfaJzRRgFP
TIqUZFog18F5lbBWC25IAU/SI/7MvPlgqcSYE6vhBPxJHxm+9+d99A1jIKJNAfTw
2iettuqPfMObbYNxjLTvNkrrt7nfrUSKUrb1fScwUogCc4Snz23f9JWcfuoZNcDt
oNYHdZUvTtFExVBS+Y9H+9oBM2GGJNM076CnjCMVxCJAmEeRZ91FqoF0ATBAPTrm
qKUWROTTq4R2vx2bINz37YF2iQ9e2oYKHJg5j0wm6Ove7LRnxRj8brbOYCSxd7Td
rW1bhHC+euMpov731oExcRtWYwtnDP6oaYePTSvC+LzlOb3KKHbvMd8251NqPAag
wEn9mOiT1Xx9Q4TrxHhwl4vdDHyRnC96fE/ZbWlSski3CcCqXgN9R1COpAL92bCl
sEnUeygfm4wbOHhC3J99p7Tgx193DzSi82JsG6C4hnJpXAUswBlcK21ULXIVah9i
J09vm6SJ2ub0zzbnF3YLyBYnohsUjazA38bBeEihhsGeczpG2g5PIfvCjCxbPPfI
zYmSVRDyqD9Yks5sCSeZpv4oi5JL7E4NY8j09ZtL4ISwzcUfws5A6beCgGVCIpEo
pZZ0/Ub00HQ/+SGasPyWjIqFh3yJIBiWlDv1Isyd2HL9s5YWIFDE2+XQDF31vesh
gZoLPqtlkSrS6LVSPfoqgvHCDFF7DI3WRq6ie7z7sdIvCf+LShzpdqRkQRLdprpb
Z+OQq6rY3surfZ/OxX+i1wI3nQxbo9stQ0qBfHtj7u6xB50uq3O8DUj6fxnmCEtm
HxEFNWpT4C1Bgkuwl2pv5hFi5z9G+9nocEkD1swQJLHY4tphS/9E4uACSgbLILUR
HKqV2xNBJ4V23IGoaU7lj/AMymPIoKR2u2nMzjoSKjJ0E9BrbGeIUW2jvIlBU9e9
hG3VwGybwb5ukrY7bVUC7k5wECj0ho/qv+e7Z+ZN5WHrLQK2ww9zP0ind8BGv8cc
Ay9vSGvlsMWtS0rxc+b7qR8rqd3j8Pq//SFldsfB8UvD+C/s1VQEIS0XTFzcFb0h
nJTwsd/nlwYX+/V3/xZozeYRiKcJRVJrvrU2Q1NBbyBl6e+lGEIFp0I+TIK+JBWw
IoRCndzD73JGP2mJPNg9maOwarX9NqSdIZor5B4l8FrODw+z5y4RHr6g0c6nDYyY
TsdD3SYP0rQb/EnoEUT0RUwo7/TNafToUhSmBdAa0Ak2eR6+tSuUBkoRjlZYTt+i
VxZymQ5MTqLEAxgzpAx5nQ1u9u+d82I+3WGdnyroDGUg8badNiVKFV3HISJt7TJN
ZblSZYRJLWrWf4UfMfZ2suJdIWQnWc/JZ7cArLpRgeW8cEu9+Z3lS7v++eefSN2f
blgDHOnWxEHeYMG6eWK8PMSs+a6vvA1I7bEovMwr+27EHH7a/UDIGDsokqTstOv9
N7cm6X9oAj3kZAFphmnPn37wwuCtpFEJ2LrL6z/MXYu/eu75vjFqizFqFjKRYI7C
Qf0REv1SUmrWZYpx8dpP9O3hVO1+Yc4yAxsYvQUGOC4ZtYWV4lYOolkEOQrHETN+
ZoLiBsJSWAPZHz1xawH5DIE3O3t1Q5vr24it01ckEWWrdiPsa7woG/5bKbXAhYke
UcNIb4OJDKAvLJ0PFT5FX8s2Kcpvcb4BVeZTsKt2guk/fpyZ2aOix5dpBxNjXJze
i78S4AS2TMOl35mDr2FI/CNpgoPhOSZdirJZ6C6zV+vLu56QxF8Y/0YP4XVmlTGN
mw8GkufQ0muugaA/ASVuYNxcMmAxCyDxuPnhHuUixwexcUofE1YMTGFq5W8NjcNR
jIYlMoXuWByZ+I1QnbXuSd2iMbO8t8WS8I7tWHoSSuGq9+GoGTnSdtjx8F3T1SnK
6bpLLlEWym48qK5cDqC6+ILk+KCkXDYCvahuxRNoFf/jfKIsvgGYo7HWJydWLJvJ
fvaazHXhfiDD6FHu/EC7VSe8xeCOF+EXOPPyLyrbhDg5fHBK2HTi9t/tmQjNRQUl
K9jHaueKXkzWGOppYjDWb+93M5pXT3UcSJkkvkZ8z1kyDCQx1x830ePCMT7ozGVL
jNbbJH+W2MPjBRtDqRr564AvAqks5mme2ynRjJX527xy0sIzcmjOfS/WCwwBtfl+
OtjNIonlBRMJ4TkROPuqoxv3X0b2QSb/ustreB11ypJRPBw4eKW6Wr/+WCskS1vb
X5/5B3exVsMtAnzXxcf18ugUo5Y1V5YKn3+mT8uJIUIjCVu+L7yHRdoK7Vt/HMSR
4mSdOVBYUrxb8hTOD5ELOCgcS16lA/ql8HjmTQdrYiNid0Ntshr5Qjk3xKhQ38jA
McxlhtsClCEeq4gusXG1aExssFIPTUPVlivTJS9fxjf6vjlPFykFJvAQ9hZHDAwG
0AwRl7xxz6SQfqjkPXhMxsVf4FW3hNVqZg3Ej444cgGcyxU9vejaexdModEAD2q8
xyFhnzl0UKG7DeXcNlMeoy2lOatQYsSsLXuSJ1TFBMvcXy/sxPlZiwF9+qo4sKQQ
50rCwQF0o73dXNxUbnXUuxUTOtjetKPIitESKMK/JO8YAQgat1dhmxOpYNs/LBRP
P1SpZAc2y3dCqDhTVs5I2wC6woZTLVlFYNIRw331C0ZgGumjQXoTJZAfRsIKWyEX
0FO5QBcAvdObFrJKuGACbAMYR3Ym8K1ejPj5mdPm4InZ18dJLAWEGQZYRvjmhm9F
tbHY3pab89+W/TT8Zvxsr83D0FVteAR0VN8jHdx84TBfAph7+29FCkj2zC7bMvgW
HQInPfZd9R/JcRltZa+DBorN4wtfoLmv4t0BnSFStWdg9jUL3Tq+weSdNdAhFLpY
MFNqHQBNAagq3aKhF/RqCsWoL02fe3upSCSPmMWOyEerqOHxqkKP2XzMmJ3TFY7u
5FKV62x11NVNh4dbkNYWGazeEP8yhP92M3PFXlNYdbYr5DPQhRiAy5nabwpnbK4y
t36Ds7P9AhCeLxmrUlamsXfLcjqInGS7gJ/TEM31KayxVoRgpFHYzbqQpK030OQL
WAQHB3JmVz4g7vxFkVhp4to/37yFmllWxJY8DJbNMEK4svPJZOgSN6UldSHTF1BL
t3+5of5DmfkEBJu2V4Brw0mKqZYirDzzyeh2E5O3f7aEWTFi3jQRObRUAR89Jz1/
Da6jOvT5Vc06CqoKFWjPiX7N+zCKt3gM7ecGs02cAUowFzbCDERpUCyH3wNSKP5E
l49/99CuBREmfg+pZmWhaPsiZH+QZmlcgGnqXP0Z2RXCqTZ5tvCCZezrGiA6BnSK
rbm8Ct5L9AcTrPmj5mlvxL/Wu7mnttegAuBZ1q/p6Tcr/s4VZbbchsb5gxCaUiOS
GVAPhBgitmG15fHHkWz2qwcjcYsiDreE5HznlDsCPiBt1WE3Hzl+yZQZAy3i3Jyz
kmpGeq6rByE6Ck+LgWQxMjQGt9tYNF03ZnFhqQt/qS3FPOmCpJuzEEQTuSTOCaBz
bbbN5bFgcRJAtl5CIGlF75dGY/yjeF2lTu7fo4zdQJ9ehmO3jd0y8DeqviYUVtct
0RKzKm22mVYNHIpjh+b4aBTVYnT73IIJ5K1EtlIb3unmO8XnGs47cqRwHAxis6dF
caY/iMN1vD/AsYExvjwK8URRGaSQsok6cKI7AZ6mknVGKMolQujVYX8ZNISD/JUB
DzLGN2kHiFEZmZmdGO+l17qQoek9QF+z+8UCf5Y7EM4CcVMmxYaLIMU91TlJ4rAS
BqyEznZslVsQ25BbqPEDUmtQzrfXoKEfy6kmMCRASOsjRHNv21AR410S5KJ+tLhs
mE9hewW15IbgIBZtbPcxemHcBIoPKk4XWrqlHJ1B2oUffNhtSxZU6afhMrz+Fv82
XqYebZcrZKLPxWkohMUVc+fBGzC8lsKQbzC3ksjGMyanpQNxlU5R0TXX4o2eJany
3XW1T/623/StDYmeMra2jw5EZIa/ZyevH5xbLadtFsHdh6gHRhMVuX49lPZHMVkO
CJd4Gi3e5XYiFE5gRHVhkWtv0b7diopIhfA2bAuKjmk0scg0RKE06Qj5/n8qTqxy
GnKYizGWt6XsGjn5qrT6FIYGG+I9ZgBIDTB+78z5qFuKmsJj91ORvQpVv1Va6BYT
wTnWRzLB7ZYhOU8sLxhD1tHLrIMF/uqxKEBmn57jGClme+1Xsw2vrJjc8Poq4QPa
Ey01A4w4ozQJ6nA7QpKUTCYtdIsCArUMkG2E1ulhQxiQc02c0DYIUbETx0dP7uch
LNfdgK3ijL45eC41DfkdrmkFEhPOOyIrFD+2LTxVDto2Wor7tSu6VnSoozRNznK0
e7hJgYcGQmqMLPRT2c5AKvvoMGmE6daEj2zyfaFr0DwDj2NAZcmW0Sx2DwjRUC15
5kjwl5FwXDbQ82UsxVtCQDkKJKdTmVm+D1YrPDcZqwr3ZWn1w6ZGcvxxg0otjIK5
wrGG9AFkNlhorHnR+YSDWFvLUscnXSxTocGbksRKtwYLujPPG/gJqRNoO82yb8ZV
G01Bqve85qs/UULI+/VmkyhJvdvKaxaiL2vpbC4qIi01zSBhUnew1o8cVWAAwgaq
orrS35+EfC5t65cbr5/1ZeKn2CcinkEQsjKmFQaSD/rXFrY7qTke+zCzsvICG5NV
XNBlW9DqNlXmSeuukknf/nTGXdx7VQaps2tmpN3uVVdjRpFY7kUzrltwH2qq363F
intTPmXnOfALiFsvUAgUESR2308Ei06jsx75PZNQNhrtDqK95EIpVImLZiqtNNGU
YJrGRfMret4oLiBCzA6a1F6bT6R292R36P5nqCKHvkrK+Id7kDWpKRMrsE8ggQTL
lFXkmzeHY2gfM8qiIctwC6Rebro2ktXjsDlg/IwjIuVuT2XstoZiqeZp2XH1jZ4R
aqMw/9mfO9RJaGAI9DiXElvcAlCt3S63wJJimRsQW4b6qciVczjH8zVUQYpgnPAT
WOvtCdfwRSjziFVRCLILsB396mvQR/dFF6L96BylcS5oiHhz46Kd6MVwxUSQCpdM
lt3oyiRzTfayuJXCj7uiK5vTLN2Ba+mGDFA6qM8XO3cOHtViRQDkyEN0sNSv/lI6
Di3Y2VWCo4UIUATBiSVU7IZ3Ep4jk8HN+hYD8Kk/LdyCnvDwZxG9LNsiYZRzMth9
UY04fX+BW75y46/SCAvLaMlABOvdBLWbGNn+qGw9sLv7OqeaPesThG056p+xVe3K
0iIsvwRyly9YvtCp3I8S9O8FX03JdeHizJukBmCCMRe0cdurV0JYomm4+hEtMn1o
chy25klhIpLyrqQfT/OC1rrn++cQkE7CMhiDjBWqWT40WX6dp9je02rO6hMkLK2T
kiO8NBZeXKoEq+4p0nGsH+e7xV/uULkdUlHewRKNYol3mqbcOhKuFj+R+P6JBrH6
nGyvPxX71DBOOVscT58tFXL5yJ8xjP1LIZE0GrvIUXTfpYZxvOacMlXjPQMFNcfr
UhrkOBAEt1NIUdxN8PmkZNW6xMLetWnC8nMLRM/EHtij4dnx46rg0nhLQcfHw52x
iZ3VUR+EIj+pOZAhzMhgJmNH2gyPktHKisruxHo5ShMvNcNK+aS5HasnvMgXqzLx
mJZAIvq2TbM7uMpzF7djUyt6LhHN0f761GDYwW340wcVKWOxSj9nAhgV25G0Ydos
UEtoknikhf4aOYzGZoCjghMTfcJVRMG18D3xXtF58l/MD5hIkQf2aaW8oYd4Vyv6
KJ2VzaM+hDz1QuBcyjsAkr+rwilUWoxTmF1AXLAdEWJnADFAegeTaHn8Np7U5VmY
1FO/PiSf9RQvwdJb+pk4tx0AcMTSSErQ574gB1cNbMmdQYbE7qnJAn/1ihgs3AvP
qW7UmZO5peFQeH+z4N3dpTrD53CrfZ5r4Cuvwd7z8xT8ipxHVkrA8dg8JQ4dkeb6
jzARmUdQOrYeh+24D3xGaH7GdGsHvW4HSQ4kaMrSWViIgjnSbPYSFAD9S8zoHOna
d7z6vn+PI4nhPnwC0e92cKeUQAMnUCWjGFFVQA0RXF2YOZa3XMbXzl9v0Pp20nwH
NsjhRlvmvbOfnZZIb0qBurQGe9kVdaGT2IHnSGqkm5IZcRaovcd0pv6+W2tbFZsM
GmxMJIoRk8RoxJfroA0W1xFP58i06ApRGm68gNDKZiboF+EKo6TGsszYw5OBbIuS
RlmRUCyymfEqO+wvNIthr3BUE+f139cwaLzMoHrH1MCLG8YW3OnunlF+tB7K80xI
Dasyl6L6b6O9Vl/MF6HzjCQn4cgXbhbSsCxkI7J4zH151W06AmQl8+BJDcceWKP6
qbdBi2cRXLLmfb3EIfuDefeVD6VvAPojo5jfTRzeWJ+XPxGBJ3xav7IUexmbAPtS
pMwnJAK7bT8Fv/gw8ZnAvtuCGK36g+xmkBXAEfbRe4MzjW6Sw4UZz9sBdeOIF70n
Pb5rw0Tlk567xU7Y0NzCJj5EEJu5qOeco0nIzMg7YI/2hJHdVs+BwuEQjiXmeMwl
poqYrY/K76+cS9H4Z8PMJ1cwArjbbuG3ibHJbFDsOeMKEXq7itP72SZ3TQfHoaoQ
c3MtoAVh8xd68B61ZdTuahflCfhukEUS8Hbz+1GaEsL1GDLp5w4hgHItCrAzqoGR
DjHsXzWEqW8xmtVnyWgOnQulbOk2+jHFhTIRDe8LZMFhq+LQQ9bPrFaIpey4FX6T
aVtI3AVRcYb73sxcc4x+Xh3ij42phiwyUXsEDx+louRc1VJzYnufbTq7ZViW8+in
+e6kbjyO8TE3LgxuCHCF+Oqq1+quc0YQHnC8tMepq2SELViXODfIYWlpMJlsvdwL
17OcGCGdeioHq0uPzcPZSRSi5nNLcOixgjEXPV4fu/CAxWqZWaczGdvm1p9wnT1G
VebRMlQVo+SOZDWseETB5xd/qvI+tTKntCYno7q4vCA0mcQz9M/QcS4hMvtYiww6
kLjffRftcRG0v43UknfAyI+6/KicVDfEy5NC2Wq+xhnXdfKBVAwH/HDymc8/FM+X
cXrO8qymgZP1jYAK1fR7heFRXTC0Too//lJNp1qK17FluSlRtO68NhmQOr60ni0e
AvhIQDrY/3AONbF/JNbUXX680ZM6IDWVUTG88+XcjrXAKv4XBPHmD4Rbqe3jA9vx
8pj8HERpp5mmoKatVtT6F3AE7JVtfUQlHURRP4lLzvjm3e8Bijdl/c00AzzgMF91
G1qa+CHfKHJbXOYB4jMG0HVBKgpYLUpWG0872bxadvNdGuRbVBQkJ5kIRUrl1pZd
C3PpKZikOn6OX76+ZZLkxRbjxNfKPkaQZzMVInEgsjqV693ONdMZSMii+DmNzjYJ
sXkw3VMHdoGzaLXJg5S2ZuGqY1VaDzDXmBEhYSAKm189j8Nikz8rh5a+jqR5e4qu
eCQkJ5E0wXQsfX+C7rEssByOWB94ltmDnBQoRAiAMiGxBc0SiXhFsDYVpGHY1X7S
wFPINQANtAT8NLodgObZx4zuO8CVdDTJOnTrDMOZcUE2dZ+Cmcm/XSUmxYGc7xP2
mVnUZ5xfJ/4m5HvRQ1Wx41vTNngnVeT3dOapcHNWDf4MqhL5vUsPtgayBQVHQbO+
5tHlQvTgnUbeTVScoNcB11NjveNkf2mhQPbQyIWwQyXYQtKrCE32Foi/qzrqfLVk
DG/6Ok4QcG2aJp3z6Mk0AQZ574jVQ6fbo8rOOYNGNTfJQ/dRu+Gigno5tkLQaBbb
WjWcu3esfSJME6IAHfzn9sTPKEca32NdSYnyaCp2kOzz7pg7ibT95yRn4Ef8npaa
ElsBcPU7OJ9KpXnx8nMj8vxBBI++Asa8OlThLAxvFA9bDXaUi2elJiK8614ebSjt
KLxV8ZlAqHuzmquwubwp/oaAuyWgCkndfGu38JX06rRmnlZ3xOtndcbw99ekDM9M
GqeXxRo8s+dgskx/FCzWp/tjJS9k82G/zJ15IIqh+eTpLqGQq9fDNiy6Te8tjumh
jiDNMXZ/g+7+TqRt1dxA2HsrRQzvKfmyTEV9DoEzWDYhdgyAIO6erXpYBz7UGrhl
2UeB+VXhqHrr/4jiKVowi6iFEJR3MVfhZYPxBaNxZriGjVkMGYWsOJ19Tl2wKwSg
0Hg7mfN6XOz/iCOLyQL8cHHSQorE4PhjnuZnSXwkpFu8R9OH2H3ToH74zXVt6OgI
8KuoKgG7zcEW0DgGBb0sWeJOLLaTcKBmSCw09ftYibfNMcdQ2cYT8mAN+JHEikGo
oogfyZn9JcXQYwh1fdVY9Kq0XuC1WzTX7QoWrCwZ8CY13J8z/O3cZ4YS0mjwx0sA
H48aWbEz2ihW9ES2I/fB6lRVIBzooYP3bcaZlzMAEXtDVUF89/25n4mXQYzfsZXR
NFvLz9wzTehzNkPt0Gz2AffqmEqLKOyLWcXyPEKRFEQe60znA6Fh8pwX7ky3QHQC
7+lNH9aWTDZZhqJh1lQcwp4AjkXfjrVq68+bDHqi2BDUV0XOFmL881+/QJKU79Yp
q8RLJhGuhwf+g7mBu51nnR4lM2f+dkWwXBabjRxopFjtsHzyw98I8VnGT6RUckcj
Xqlr/V4M9sBk2z/GcXl4tUj6gYmu08a4c4xBWdWPd0EhRap85rtbvibQAoKFJ9Gc
tYzF8apGAdbCEzWT/AuKeDJcBmsAGD/GMTdXkYsq1QvCBzmWBK6HnwmJEGg4uNzt
jYBEto8PZjK5oh6wFC5EswSeeta3dZhYGWVO8l3U9onWLInLuSGSDsFboJB9SuJq
k2noLsAFZunCrLwM1acHw8lWzdhpFgE6lBJ9hpQhR/H9AhV73Qu6b3aseBCdY0WX
A8dKKQrnjM4Qfn6NxHOpevXyc3KzzKR6WXHkieZ2dkFKWyOKLIbyCpDTC8CkqnCh
+h5bWjB8Ax8ucXHXgr8zLn+SKAwjB+7hlKHX6JE9baDkWlUCOj/PAxGRL4GZlkIx
8qTJjR3oRz7DeS7B8J1EnqBd4EfoR8GmPIl8Jrm5/rf//8MVtgSjFh5N0K7XXJWM
Xbn2o4LFhXQluKNGyQLDl4addTuluBHniONI27i4HtxWvOMfAOISoM54WK0eNTpM
x0UVi+OhghKi7IM4mL+xUomvtPG36RsyBC1L0NruphToXG+DP31Ya6T1zeNLIc0R
jdZXhgFiqrGwUf0w0tTOkQWje6QnqyqnDFQ1lXAz5V/RFBB82uosXP83/7ckFq8J
MGhzvLnBJa+FLgoDyPOCQMLoZl/KPdDZ9MPPNDwSLYulZsn7so5VCnPNIHeXfeby
StUuJPOk/iMQzrM1yOSojvkudfJQ1EGW3tp8uaVoESsmKQtSKB8QdNopNF8RyHVj
7NltrvBMVsB9apYW2uGjhRRNg8n6iAE9ejRfm2uXDPduJVbzMgBa/K3gPIeExiXF
L+U/zMOwWYZiU2cDQzCMdAfP/uNBr5pY8qowkBQp/Qlx5AyvKZHGLyMIGh3igZie
oI4zYR4LY31DHlhrG5x+7sCaJJgnfxOhsVmrPu0upfOomPbDnAyCZHzrPAUt9uX6
OBgnNogbxNBkElKUGQdOuHcsJ9z5F4dYfD5ZtS9uv/2Dg6q9sCVUcSiiMm0sF66r
E4kEYku0YoFRgE0Y3o5QMCZINRvSkx8mPjGw2Jt1Dss5xNGrkU6ZWu92BneRa6dM
35+wvguqxllE0Ne0rdeWYNJwRVO2mcYYBmVTw+BxtWXDISMylJR8citNEXlpDYjf
F74Eutq6aTtSq4h39fN24pdw3rRL02tFfiU6RmFzsXwhsGdLh01lzvQyScnVkL1V
xVysyFOXgrp0sppZzAP7cWtx17izuQwOiqsIGJf8LpxZut+6NSvKTY+uhfSS1W+X
gnw88TkFJRg1sDGOCDVRsLmCbAuvCE+Oz0q19YFJ9TgZxaAdJu9hIwh01T/qzAg5
C5N45EeSDWll5XcgicztE0boIoB+ebmEyrladWeVc8Cg+rohrHu/xdF+wLJ37bP8
W8NcbouZenVUcUZceLsOhOpanWePymwSkEa9AVmnQqOYjp3dP78PMlrDVjRTk+P2
DL7B6z/yP5uB6fjpCo0VSdr9zgKXCxVwyeEMSQgZ4wJg29srUmgIkJjKDuc1Oy3O
wpW718TvHfim88OqlFnkhBwbaCKdi+qb5SbF4en6bzUpFxWKtGz8yhKsJtehJQ5l
pzV543rb+2af+sQdXpjIRfYMBlVijq+qkitknorG1dbAZKnpb82CHd/uUbLO0KDM
O6ZfKM1Ehb19KwMxy96qsDHwfVrnIsUNeUi7GjnjMkbbfXCYav/2G9JMLkhZ6ywR
I6M7zfjiYgL9L/HoavYEThHSxdrg9kHWqc++ia3ngKNltum5HzlyfGfeqZUbQL6Z
hFw7S+rN55rbr8juHuxC9QnzA7fzJ9u6nd0hmBUHCKBtnfqjMd98DmvOQY82zp7K
SqpZOpyt8LUyB9sYUF/GcakTUj0RJMS7Hv+SWqMV7iOH92Hspk2euCXOYZgCl5eF
9L9cSgF+VTcwi24dKNwOCkyy7BVSUO1oJJPbxlLAZYRHTjrYXBN4jfL2mHA6BeCU
/HHrVMUuIxezl5bmIcxiyEagvMSMteVk+8Hw5mpw5+aAEWeAJn6Wc1v8tRyWrEd4
Ysig3UDH7PwH9Na8B0C/P3skXnFSGPsK5ZqMmP1GSJVLEKafI1mFMFYXb/MpIx+w
6MBuOf50eCjGr5A916C2/iuPhhKRID3D2EUdbEg4NNSuKU6L2Ai1oIPl8Z8rzZrn
JCuWYwDpDvQOORG7kTw/N5ArhxX3SXM1q4HjcujNF+7jskClcCtYsXAxu03n8dgc
bYsGXA8YVzB3dTTsD8gDCLAQyzB6RjRyEGNCCBBlt2LTEIY63uRd1aZVB7iEGsD7
ope2z/kJ3K3VTbbRBKHFEsFhNbD/2tV52FCEDplY3Ltmjh7ibLeh/nRGkhnh4eOu
UwLFabPoiiaDfw9/PbhiZCIDXWxRw5X1Kk3/zEsrqJwGS917Tg6OXF+m7oszZTbl
98XV8nM1R4NX81+3PiLt3y0KuJ+bpMixCQ3NuD5jvzyjwx65aCGEmQPmnC3KiyxZ
SL4yoaqwk3ubLdq4g5auRI+pXcbub5HkYZYS1GZSvsqWS2VBiuOlNP/y2HaHaW9h
oK022GPlvW+u4qyQcLXYHP/pbYP6P7sVfPEWpSA9klRLdO6q+XnQOIR8L7Ia2pX3
p0AR9LsBAZwbErDnKsG4XvYszHVh0DpsATbzFqcGsLgzGNwtdBDIJ/5YGMfNXMhR
iAGJ1DDM8JkYUJr1OoyJOV794Cq0njEjoo306RGbZBv649JMRlbSXNNGgJIlUCJU
aVWxokPT0amuI+0JOSGUO06NWmvrDI0RUGlDQ+9YtEI4HJvhwAr9M+GjGdRbv0xD
EM6poJO4A1opMjFpfcbPl+sr/XFcIhVmCkOGOx0QC0FOoLReUNF+qS9ECERaHGJN
8AvqROCuEf8SROzg8us6+oW/07ETs0JLaLDAuf2PBymWEPEsySnJ23jbDCPbrlCC
b0OoZRNZISs2QjidgPhDmetTqG532qbuXXIAFE2UEYNVaYAnE0kOfqQgsWfwH7uu
R06oGGt3pklw6tI78TGQftCF7lHRZP+iBcB2ypR+joAhLFk3lZvsX/PlaVWevWaJ
/GhAYqJh7remlLB1X6ARxMxcKXhWREiHz7zdgC5gguD/7Xoamafijnk23PYTMSeW
rFczVcHuKz8VwP0+mUqC7/Qu9RwbvvHmscjNGEmwhlFOvI5cfdJMfD+zTwhi4mBX
XZ925xTak6CHOc9Wg6Z4NtTTRvWgcf4ZB7TN3GmR2bmnZNw6DjYoFDp79R97kBCM
/1emMTnjvGGv9Yd0+HKWcUXHs51SYqDKY7do2Vbt6L9isjrnD9m7XCCKvmH8J8+a
fNYHKP2E+ETP4gkWZeIsbuUTa4bm2Rg6OXhH1JFNFgcmxdopocVTwhedvpQzVqGD
8hEDA3QRpa7+256QQ7EKu/4O0yn+Q8RkXC6APBIEnIKSjuenhIncamzYZqq4u03H
wBTpRcP6jqzUSmhZ7nRG7xUu5qw5C8uHLxT903yFwta2CBRghNJBpqpHKNctGUPp
8dk4xsC27414AHoa/hzuPBzq36czMn+Tb8sRs4W6sdrtl3eiIFAdsG30Y3XUaY2L
9or4ZZiU1eN4oicNgVX+G/O2uxB2haaO+qL+fWMY4BI+UVYKQob+lk0u3HU4NyhY
JkCDrVHwTZJJmdHcY/yvilKQyBvZRvj+ZQcJd8ZZSnACiO1/QNMI8VdgW8nE22e6
haxSC1BCYed0OYcbH2Z7zBQqWqxwltUv0L8T9vXnhXPn+asU90petNZrguTqCxKr
JXUeHnKZKFlqwhmRMyA0XjH8/dO3g+lPkRh0KjcSl7Bfn+blNOPiUAbiNLEOtDw5
g7zICQ6PIhw37hZLCvBgIBfpV4tZ6GhrnkwO6sZrOjilyJnVgdSTXyDSOx+v5iFg
3jgbsdtfnWjRf4dmqIOwKClkcWk3B0bAlFQaDP1JhR+qMz1UqYMMb84xOSi48YJU
wHE0W4hhUhtIUDCjnJB2zotvFuUTJZGZHdq7SyZQ6b/CtzAh4aw79mf+/m/w6hSB
f9ZDuSLwSjbjxnZqdxnJlf2n7KAUKGgHisv2Thyg1zXilsVqdkgCAwIkGSwpXiVn
58MDVrvRfAhKUbAP8G+hZqQ8BB9basyvaHa5eXsma/qO7aH+147y9p3A8yUEiO7u
cdqxQGMaQUp8lAl/Vyk/e8N/oIcFriA2V/Ms2VxkjfeKwtB7RFb84Oq9R2J/Mzmp
pPrKtzl1y/O41uQp0Hstq8YQB/3o5gem74dzkLzwLjz8S2az20FtZI/IFXwISkvL
82/IMCahBgTrxAs5BUAQV7wj731AuzzM1le8fRgn5AxHccpKibrm41FHXWLOUlGQ
Y/ce59cxtBR2qGg5CCkVgLcUuGUdJ4hPjKQXb1zylHnH3bI8Tgf0cKaeltRAAFqB
5bUTNup+zSt6FCjPQik/irJOvD7lNKQDBfnIJ40bUR8WIx86qOOTR19BLcc0Nv6U
FVjjbpwk4i/uD30Gx+gSnGRD4C7WRktWpV+HHL/fO07VoXw9+QxFRG2Pjpz4e6ab
kP6zI2McWSd8k5YtEjxm9B8gs7WhkfdqgLiwgpQ4JtdsGa0AXTxYSo7Ts5aVdzTO
5hfn+yxovB+jC25CQRnrv4RDu9aVzWjYKqUd5q4S3zvP4vnOJlvEzi01/JWfuyK0
9tL4rHwSfKYCyVYLnTlP2h2Y0ZsPvhSMDcX4saGOhp2gGii3zm8MDY0kH1VBeeCW
iDoyX+qPRweb1x/AcTqm31s2OV3iACCv0CPKtbaXD1uB+qF2HslS+/f9ckPUED7F
Et8OiDyiyb4y/t9sdKkGJUM5ROLc3yQNvHVdeRbdgcIFqj6cnt6oeyPzo/2mUXKc
piSQap3tVTMGpNCzpAOfkjC03xxnSayJKVrr+PzajiFL1h+7oa0Irzm4X2292VdQ
F6IwWTbo1M3dtdNXzYceL5NfpLR5oOOMbBcWc2CFyDVNy9cvdw9Uv/Fz6YiGWVtN
VFXv66Cu2dBkfVNOLa6KmANvu0R6QtamanjwG7VKmMzBTHbtzImMNRnHHvUMSg7w
e8gHhS5jFrLxq6xeu0PKslPhVJypBL8XRZPwCSaxwXHR1swUWMYZv070U6wzF4/a
opWeyCc9BpNGB09Dn183vATTsISCeP3MagwWp6zK9hrNBmoMRcVbUOxUVEhPoJvq
txIyCiQ9PyUPGkvLXoVjNkRBTwh5yC6L3enbFrWihZqAALSE/5Nm5MVFiiqnCbqL
1Kr6HP/xO5GIOLtLacwrs4Dan7yei2pbeEIyi05HkJVztC3uocxyUTYXqJOLq3gB
KI2J3JwbzvsGT3MTzYwa64iW1E9cOk9Y+6sSUeFECYQFice3Za89hsN2DygNvT36
XTZ84ELs/cqPHE1hbCQn4B6ce1tNsOawEU4wRATHwu+I97kSL4PbVhb8b/rBBjgX
QYAzaZj5D3IrzsZm1f7+SHCG9MtB6p0emvmofyX9az8YGxwbbGd8wa6iwvVpSFuu
EvYhP7AwqgMiTVZlx/9jExqWA5sjvy582FMQHkqtrc1rLc0Hg7qMGOKE3j/eX7VC
Fqj9PKQy8XfvgbzJ8flRA02MDfHr7veiKK5KekC0IxBoK3ygjZBfsAAckX7KzkUI
WUymcvQmEeoU6Ylp2vVhygj4dqe6l6q2te3LmQvgmi9nQZZ7w//i0WxQxlc1bWUR
FyaqlxUoy1RZ5q9kq8aDb9kZtFH/61tmd2FquRQ/Qr4P3gWQdtrdAafd8XXjoKpS
fzYFqL34Sq6anUPc1uoYuFb8v0761jDjhUPzA4nRGGDwhtpLSGuGfLgu5luJPuTK
41i3CnOQj5plFyV7kbrdrCXpdYxgXMTScBffqamnCJAikvrJis70jMgrgOZosxJC
seR+KicxWzcubDBO2oJKjZW701pds3wpHekJpMzcPdu91/ZMkaiYLFHyEFMWHyMB
dbDMhBcT4ts6djb/VkWOqy9yYM7IiXVWFibkB6IgDvvVnX8CHiRl2LmGDBRzu6Up
EoeEr8Az6iBNoOB3O2/9Ds8bzPz14ywiyJJDvOf0n26+uK/ANcBJN1MeD+C/WV/u
dB6wMfgugst3W7CIvqCOkP2o9PzN3vHe9+E/odiSb8frAMlWUzBXRr1EMKaZXMlu
ycHxqHDkBNTisdGpscZLnO2KdOT9NQZws8lkWrONz+8Ft8dKsMFERRz3ZPugBxGi
D+JAvjD7az6ymXeu/p3xig4DzHnCT2I7GJJ6abrWBF0Prkwzhf57sAp9tx4KV9eC
GWbLhprfwetEI7jKRo8JF4JxsU/nv8son7tXlh41Tg61xXvCpO6IVm+uJ8hUmREo
qzX+yf8cPG8ORnhjPYmqhE/79h56bjEKuWh4g42kyMz+VsbEmfa0jeoJRRuen+7N
qr0X4RD+Ww6uDO9Ds6P01twJdBbcTeR8ng0aGgF0N1LoBLlUnaE1squJ8ns3HtAI
hqzlQXRl4qPNy2M7L7iwMs+pCjFjrLV5NhgTZJX+aITc8g4mFX0giwjny4et5FGd
pLR4fBQcjwELSowP30EejQMh3UKD4ru8jD2oifAeQZ5zO0/dGbadIl0HzFJU6XYG
oi+sujJoGkW7FmpDjal9ySNE0YWTs9Ec3jfZW6tuBBcxe2lwCzS+/CvjPwSYddtT
QNNG++QRbusR9H4Iv4uRysh2TIz8hTIkgVq7atidveTzDo3hiFVwWhCeKkAaqMEy
odZJaXvWaaEnH0JAl3kYHUCdziVkgAbICdR9PhzcVFRcQNl/+z5Pw/VW3SWNBcKd
8fb0gxghVpnPjvdZvlMnRJ2Xle4OaG/QSINb6F7B8S+o0f1CEyEmDrYCPIf7eX0S
XNoPgJHsAG560J6o6165ijllamYDgKHudiGByWCzYgtSY//708xVPnDW63CTk17v
StfzqXaCnbZz67ueA7JzbESOoEKQzIiH8iDpLr0vc9ktTcuqKF7XGFr2yrMO6fLK
LYxKBotTnNg+TLDohgVFgbHtPK5dfMYF2mpQwr8/rpEEFi+dXYfG2ZSYSe79aRWr
bR3J2ItQfXyxqntqbnMLCVx+kCqe68jXytp8QKmXuN34k1ovrFxsNN/vgLGUDP35
wmipW6QLYjE9QprcinSFHluY3S9j3cxfVfmMy2r8z9fPqheN5Cjj3QxsP8V67B1y
lARPnqqDn+Oq/Lm4bqJHLEfGXMba30+aBL6Z0bLtwLlUo/zOw80oyh5FgvU/tmDT
1Kyt2iMHWc6obHiCM0i0M7nqO66moe37ZezBc3awa8By/YGSanwgbd5vwifyQFKb
Qlhe4XHNjSwINVejB0FsocUDBSPu7kzH3l219HVvHEgh+Yz+KisOmNYa5x53/4gv
kZlbn2itCjfCKZ+4+LNU6aJ0q0EW2i6lZ4cgK+60HBq5ISNlA9OYW8AMY67+mLgD
Lt9bDXX3/m/GwmPXq3DxNm2yllMTY+9L/9zKuFcu0XSU8UUaVeoxlr/k0zqSPWJe
H4zKuJzSXJ1DFm2mhp+WHyBJw5RNU4w0OkkArrN2G/K/+vs5zWcPjUyaVSxyydTU
SsgZHogO3svdz/lpLHkVy0Mh+hP+RtWkkoR9vk7ACzQPbjcMBDkAMItKhL/yASQ3
i57YXmzrDIYWkFq/x3V/ewvZRZXSc/gpD3DbekB3FNvGEK8Zi+isxD7srGII1Nnf
8nBQ/Ub+/6GBUxroLPtb2VXjsmRTPB1ub0BSkezlns3ut4G1hWjWt6zQFlCjlxX5
5WdA3IXwqYbanATLgajTMR8wWA2ufscejKdnOnqIkYtuQvdRazC66Cd0bERs3oO2
qaVCN5c6JVOslXyTTloxVocWmwBq3+DdXFii/tOzHsIu9MNs2yNs3SxYt/elroPl
fAAPXO9KAYarmFFAwPVphvellwRBLu2VNhyiW4FMLPCW1E1C7ur7TewkBxPW47JG
gWUl2+CJFvOLqVt5zKhjuy97UmUdowxml6ELXIsEnfaVYqi8QoOuddmRyjR0cZi2
qfa2ubeiyZkU+NuTFWwJQR4v+X4HlOeW0pgcYcOxh6RXSoluKNxY8qP47yhgZEpG
X63DiRuhn9haDIOR/FCUJGHM52dsgkkKg0vGMXfvmX9c4LC12hItub9G4awIbPJb
TSeV416fYCTzuWUYCdOat/ZwjODHl5y492DWSek5q6shU8i2a92aahwHfFOr60qt
NmME67l0NVLtyGeMq+aCTOZWORJ64Y63pKnxV503YEOq42YKsZNdnqDqz8/y0yU8
yYmEtzVAoj4WgOH6p2rggV6O474eHiTlQS3GeQjCKq+bZiFsCHEqZe6I0rgB9dKH
dWXXjL2RAwtdz5KlVdsQ6zl6bz0ze36h0x+vw9jvg334fh+sEfGxNeor/Rfmrsc+
SNIuUw4W1QGEa4bUhLkksFCIbKaXkFMGspAdRxD1YEHAB0FyetEykZ7MDMXq9Ia9
4p3g+7ZblwimH2HwJat6rC192iZJeqel3xKiq9W5/Wv8z1n6rygjJ5Tm7EVXrdUf
QG5rGz//EaJiYjRHufLX/N6gHX/TY7IrqXyUYNfGxKzQT0yMUpQqtJck9UQPcECl
pZJiElt2hfJF9kdtTIFnDR+AIyhF9wWFibKTTPKgQL9h0c86cEpJiIUQTYi3Q7Mk
QVpsOeu7kATBbsxToLuvAe7xqCZDh2CgimmTYa/5nW+zlz0+OlfQl7CAmLZO9HOp
c5nS+vhIEl6Do6BHF9yH7NOdYP2ZrvLXCeO/luYXN2+jgoFOZtzZXlqasZ8DeUNi
Y/frgJFH7HeyQEfuvnpg26jhW06pxUrOlbB/IjcnSeSWVJT6hoxSMf/r+apyQXxQ
IyA8hKud8i7YEijF0DgywXXsgasHS8hgz0HyW4vP6o3PqUWkaL2/v2RaU8OX26LW
/xATmhClA/NnfY1UTBjqNCAioRuFXj4VFqIkIXY4UVI9SKVgTysg8swbzv80bxvw
BOHclxx0/ICrqa9Eoroj5/t71qhjNdEw2PweW2xITJ8yHgo4RIyVcdEqB/jYTazg
Xr584jKHhw9UvSe/9TKoDqnJHChidQaNIbfLznLx9cG/5CDlBy8gmht8ksZMPRPu
ojz3jrJq5xnlLgUNSsH/frIa8cu5dcRxcomRBAsepS47Lok+xvCc+hEg/FQpFg4p
MsNFxBPWaNcBARO2l4fyLu8A0F0PEn1NiYmjFILMR6C5kyHhvHgLEmZup6hA+1/c
PE8gVo9NTjalVXnb4wZJFgWw9EUd/ejOdIxyRAAK86r5lFPOaThm/+EAR1Xbmy0D
fGXC2aMnwo3xKlhkf7sBKx3Ykv2+obWfnQndgI5o14J01CqkE4eTHkk0aSrKTLlM
7OA1+nCU1FrzdQpGxkEA5GQthT/bZAbwY6wEKZ0fFJ9A5nMxpEDpFA5BGbKYZVxR
qcLRAStqTnqdVMmbGyGFhDUJMH2UuOV4SNQLkcvYLZ513CRJWQ6fgT5rOvvBDmcS
05t3RpyA3n/kNIUer4ucxZ9QSuFloQKRYXsMS6aMEcc2wngnq7xKNjWQaOPaABRw
zTmnWDCIWA8rRresyUUnTqW8/6OElIBdPQ8AW1gcPmRi1Y2PJyXfT4BBU+X9OmCT
cFC17v5Ihi1s2QKMxBkxJYthT8bgr/oiXJ9SBfUpviA1oO8bFkCTZLntrxvG7Bq6
OG/6R/hajYZKxq8Ajm5ai4IrVD3gHF1Lf68hzQ0znkudqcsVXxwB85XL0hqcP6Dp
mp+Qs5vB9jX+fdBgv7lJAMD0RIBqb0ERpxBE/JfeI99D3Xc0f9COXmRHWRRwxe5P
SRs33b/EQ0YlnSc+2CVsFZfhZZwc1lYlWmApGOvPWOPup4wlTZWf7olPCoRTBTA6
+uPjKOneJme4ynRgOxWLw3hNQv6jkJVJDZvNVHjJ2+7Ovqco7ETA/Ji5R3z2LjcE
Qt/nAgZWO3ALXMtSbCagaDxMIhBSTLv3ElSvgR7XIYHU3TcmzJL8BY28chtR0mko
bK1+NIJtQm3k1cU53Xp7aNOQOJquL8ZK5JnH7ienpgCEPOkz1/SZwN03RHeGy7I2
e4vgSoFQptdelJ13OHY9PW7KW/A1yi2KXW8TJMnoJC5E8/8V2OPOgNLEHQ8+8xi4
K+0L8pBCdLTJ+lyKsYKa1rvE311zyZY60lCZ1x4m6FuBmhbfOyZWCtQaNZYM5HI6
FgrI92aVm+nc/Ubr8Dh5qAy8HND8doKEyMZegZeG0mfUpXd6Cqbup9ouhL0EDn1E
ATd3bSjbv0LTS5fA0E6t+Z0rbdbafc8ySTa1iJpr37nHWiELfJBCybqQct2p9R4k
ti1MtOu6Osgz3mr0ie+AT0RftrMq1jSS+tLI7/qS7z/+ycea7YpUjCIUaY4GYHog
Kz5O8+B0Ihv4Ja2gnyYYNjbU238LSNnoOBF2xtN9dscscDIBkE/QVsB8Xwo3NNWT
qK9v18sOACoFvhOcerNX0ZX9kjkamiB6VwxhURXDJbIngjf9iTInahfdwGMqMqI0
u+o4PiNlbzVMIkPywOyGjJsGrmZJPgtVlgDOaF4MOi8aeXGQkp9haQsMgonp4I0G
GIAzayjecP56pXMTQhU8fmDQJGStF5qpOrvmCr8Dw7iV1bdS6eCQKgnM8EKsPVyX
tH4Ks/WARCUcBHar9d/AD2MuTKC+BfVEObMgk89PydkwguZXGm78Zl84rhacBGai
MkIz+0dwcgSqfrUwjIA5ldFGcojOwJGlQCiP/HFdq7wNe5h3Y7yvEW3QDPNGxmlg
a6BBZWeEfFNCjEyG1WvWwzV3++X1bJBqWvz1ijEAKi7LicGhOQkySqo169yGOk0V
zwuqHG4H4PE3mrfDAUNnp8px96JV+8ZIdG4RH4KPtAKpJG7Gbx216COtWleMwN84
mHFC+K9IyQJgFMxzVR7to6HD8R8rP3BUMAYJ+3k89yI60NkZBIP3k4m+c+GR57+4
gTcwYUwFn3C1pdtYQfSGGyAwfaL1AJVUGzSX9pYN5TxTA/D8eF7s4QlgnRxqD9pp
mIfdLNGrELXcg3iyQ+PKtq/EO+3XnxD/+4730R/WcD8D7ercVwRvAHXLy6IxcWrB
smLOqfkzgh8+qCT4RiVnC/wg+3GsUwhpwqlV5AWus+H3g1JCfBJEelb2M+IBl056
w9HIn301sorJ02TNzWIJnIyO1ck0IIwcEVIHKFjVBFHesxUsmMpTRKXJ4xPKtBwr
ZjkeAxTg4bYFWr/W95GazxZVac5qBF2q4yZ0WiGd20ek9t1VV/GcakZqloep/G5X
6/OJGhyInAevAq/HG634nYda2L4hX+X0hvyTrgtzWFkHCAizh7MmBzMMG1bwZUqJ
ukxKiighNzOmgWT4QzGaG5ENuFS/Byb2yATcSix4fcBkZk76jee/Gt5y9tqoqNU2
qoLQlrsxbF0E67NpjacKe1GUaLuSQsk7eCt5tURKWxymRc5qrXL8tmA86SyGZWIZ
B6/rgtbchBq5G0AjtJHqtf+bhyDTiAFqsUpNMqTsvK3NG5LLaXgWo2z4FCXRZWWG
MBVq7f1xw7r+4gEsfHki9zYzb2Wx2rdOjvPhyNGjButoff3nhRi/JL2VKYZiQT6R
qTUQdymJkaCxSSGyV7TR8TR0BCPUvO5Cu+/17p24jmSycSC58oriVaybajddrAub
+6AXzGSnAFFHFDEhluJyCeg8vlhK6Yj+ADUD2dQa8aYPxFShKVJAQa06JfobQs6H
iLL2AZAGQrtm3Zjij1rA1hiIHFmoykz/8JAaY5vKW/qOq2PJgI4QV4VNlx0uKNTr
T5WOsfRWMt0EC84dx3qlOSgdzdx82oc2CcwQIdvY8f+Fx2L1mWuP+XtJPytjBIxo
UlLl1fkKUyfGJmjpIq1QaluixZ+8ILhliAWTWzRUZZajgyIWFlx0nPLG2M8ItqJ/
33ARPjq//hUVFIzFBy7eoJFhYPqBDMe3KiDXQ5FIlk6odqUxihh4+BvgXCYpyeIm
oVFJoCMaPiJ9EF6gVsVKNFuYvRN6KhZyJGKMUwOh/CkuM4JrBbrQHZcsTjEuxVNI
qevMRR5OsU2cEBeND9eG5RVBbIQxuV4fnMiuXk9mINfYywI12UHotGEgMlkl+8Zi
BVJhnAqqa+HzvF0M+1sMBDXBFODg0YKlt4vMAukQLoIsBG0mulchMOcDKoQUst7g
xLEAfME1sC0aqicecJ47sx6075kY2e2vVgU289Q4ayzLRoEcNmx85Pg8cGNEVJgS
3A9GwRAhaJzcwQcEMcb6i9Bt9EIa4P1NU+ksuqsNYiAdJLxOvXWe6PjvxrtiXocY
ejD9lfhiq2avpH0nnxAp9RIanXhQbzwmijJWDnAjBqoBW5z8ePCXAlyIFndjptmT
Kp4+6XJdaIVHxZBtLJ6VmGypfURR5B+q8jAJIpO0pzDWXEZUiMR9tR4J7vKHJjuJ
zmfT4IKUlzAk5H4sSymMKErhsR2eIfGqPokCX8rjaJQV0QFJvz3DPmgo8hxcAL0a
xQCEdqD5SxCEEEEls8GpJL91TnJjpRk8WhaOq/KikfW7Kftf//I5PJvbf62rCZE+
rNtve7tyjkZA9ekFKT4HfY4KEyGM/5DjOGvT6a21Mw8E+KNeZPCQ/v+Sg0kmCqZN
7OoQiZi43tkdTDocptHHot3wi1JCipyMl4NqNbQbUJAUMzMqGNOn7px/KMm0CiRA
v4AbaIDy0iZ0+1zluHPm1c6FTaA3aefy2LIslZvveirP3b3yqdscO/XbqFUemI1d
TYkvnI8ZmnmxYlpscS9bezSvmp2e5izfx1JPfJ51JFHcI8B/rwlBcSA18SEaKNeM
b2lBGRT2c3Hi9R3iMKPH9yhe7yakCEOuahdI9WSeHrzrKjq4Nqz9rzDyT68zvL5Z
QzBFfR0NjPz8wV/+uNq1aTsd5WcXGiHEBUntyVYNpEd9plizSeT0KSUhYIM0XqIY
dgxBefDZ7A3t7vhHYMtlHxlbq+iY3uIf19henYXgGY3LLfz1PMJo9A9rCre6vKIU
/5N5jKNTZp1UosUmCmFPUYCtgbb/aIjnpV+ct6zK7/hdHW37vB5X9cVZBP0dLM1Z
rYFHHT5rOWw05Rtrs+k5q/vcjulZDukYedRcJJygFGvfv7SmPfz44H6s11PRjZVo
96ZjuPyr5n0tlnMih9I6nEpiklLNQfbAfsP88p2tpw2EKdQDnieYq3HLsrLqVACV
EW0gbrryd3V8QTTxTK41FRHWCrNLT0c3JbRQq6CQoSqqESz2qevBrbWhyrddWiY5
r+fcT7DIxC7emkk2ahEmk1GyG35upZ0b5LUJx+BQBjTnoBdQiEIcMqsD3wXB0YFo
Ik4SKk3OraP0Hnv5rPtdnrLB5MtKGwbcynhQZXIP5r/1gZTJI9l6RCmflPSiF8gm
ooGBNup/bfcSkFz0r/9B9+7b9OPTJJMXzhtdZtSgEohdnD6cNID4iLmIE/lmukb+
zCip1m8/OUnJk5l3z18eb5Esp0iEeCsM/p655V3PPmt5UCE5CHLWVbd3qP4Hixfq
hvGRKpOBBvxMQ8WmcrWvgEdTS4T9ZKi1WxJtD0pj9KxbNa6PakiAVa/QlSf71T4+
yMtG8jPzqR0TRkOkjRityKm18v6MV5x3AbN+zxuvczfHmiZeqz3TYPUw1WK71gUK
7QCYecY4l3YBu8Ml4c4xeVzrTPltSKRpFSgEP3FwG2ooKg3HpuqsjRKfa3FDVvsF
gu5VI88utAjTrHtrXCcHCrll+SKTmhl7ld7CF5RHwuwZfYyIm1g2nHWmhzRWNVDx
kFWW7HBToLhAAGAuMOBlbr4MMv4XwZMhMVyM3R8viRHQdWN8ODxRyfJAzeplL893
aRLDY+zcfajULN8MBk8iadnQTNg6KzZl1Yoxai24IbiKK2DhqcaDU7GvdspwHswL
krbD4vWeQvbQCsN1h5XLU2YHBJ0mWHEa0nihrB1DWR9sPlevTTfd76KyMgFNB1DM
GsqBJ2n4qyX1/gwkuGysPZsOenh/kiUKrxd8LXVQ+YB0QGR9ZPY0Nqf2yX47yIjr
PbnHEGx/ufK/2BLLBB18YDY620KWb+Zvang6d+5y1TrpB9BdxeUJiQH2hky/G0kK
+1zOsW1DblVmEq1BOP/samXk+gADB3q0P2FcouAoZ+KynqhpUyn/IudyYfcoNMIr
KZ0IJ7F8bibr5dE2J+BpQGInMOeI8ESikURR/ZiTQrlW/3MVXvLfFcbEr0FOeauV
4Bs5YXzZ68Mt2uAInKlXaBoOp+QfHznu6WClwWMfce/CM0tnTyPD5TTjy9uK5FpC
dBxwRBiOjyKVGWQ7omVGKxLVSDf11wXVbyQVUt9PNbXbBNS5PD/MXPUpurDGa8KZ
TYLq/9vlmsWoLH4QWwv2d6D0I5Ju9TTOQcRzYBXa6kmCqxQpdR+mnrHSE2N6GqOO
Ao42hKMr0D4CbfvApLxgIIxXIUMKfM3PF6joQtC/RlHxa5feJCPQTDrrOvBvAH0r
NvF5vIiHRAkRrcgzU7zb7F4vShNaCJ46hS3uyI8VDikfTQvjatMTsLUU0TunnlmM
JuwuQxZFBDWBoWsBCl4VfvPJrqtZlwaAhFTwNfMstSoKeFNpWtQL0KWrGiKYthXR
c7b5OCPWSnjE+E2gmglFdx4expXOIWk4Vn4b+7KJ5becaoxsyY07PRa/aQce/X9i
2+bkWMbxcnYwo8F9ml58ug7WXvrRBnKem0nG/9Ei+vCU3JaArio0wNXe7jxRhMUT
wwiyslOsWI2dRIB7F/STfyIU6sXTzAc1BHKT6N1ZHG7IMORSET7w4hLfq9HouTdU
4dba2LovTCI39MZPGxSjM7pOxP36+YtGB8pfltRkMyEbNOyQ5GxYwjGrsF0Rw3EZ
sRgX0MQyPk8EAIm1CZpmy84lmvjOViSxK81ur+A5tl0/3yV+9fyVtwNIxcslHaEZ
r5MCisYnSsZ5LmOdaPsI34woSK5qJJg8o3598UY2cVsT7xT2LPs4+qrNWlqJsHbn
0QH5YvOFwTSG1KK+ZYRCs6vrTCnEf9E7cASn5b1VFKg6/lcuswY0kKktoWhYCGET
3O3kNWilU+ZGXT66gAicKKGMt684vQeWfQdfD+BzC+gNkZ1CmC2KJb7AetqWkEDK
Ru3pBN4twTH/LVDIY9xDgxA1nrpRXZ9SIsTynqQBKIdjd7so+NVGqyrNi7RHrp0G
DwWY+GXNYWjNVGYxsRkeOz8dD5c8xotwnAzn15qMMMemK3PruwPfKxDAMUUyewEQ
6Bcr+ss9jWqfV5TZmCi01M8jo3FO69FLOJP9wHXgJvcg831xe3E2frYx43H1LuPg
JGqZrqGjKCxzR913RMaRPuv6CGkYsEfSd9/37gObEojxrLsG/tUPvYDhFA6iZKOd
7G9XdXa4IR0Dgmg6d6xGmSrVHhULU975oqllRKwxp66aynMyLkgsnHSWMb97GSY2
trKkFeILGyfAcR3Ur6S3F7SZx+qloNyK9BxkR2YjOF77c3m6S5jTR9uegBkfFrED
CtJUTV7lEdgq/TgqQf3IHoM7q2mM5jJbmMufWZaE1DZxXElm29I4rjcKJMhZgdWj
GH/lwxeb8F6pUnWSPs1W44Lq6fsEptuullwYl43knPR3mfvQsrFKZNXBZYsmgAi5
8xvQy6SLHLHAmWnfY/7djIrUWssAQek9GbYxTXGZ+RCYX2OVaHGTKhglFNdZR2Jj
JFffz5lUa9f8ByC6VQlQ9qwPvfq05qadTGEwXotbE4D2y1eTFiKPWkFwhRWMkUsH
ibx3ddu7nOesoj04YIbbafbpaJ90k3xdEzetuCP38NttHcdaAmvK4aSY3PaKh4dv
/nZVjG+AO7gmrZkN5aoam+ap0h29C2NzS8ZfJvrNnZ7NE7ZkyCLlHIopb1B3p8to
4pNAATd0lB6vs248ciTQax/o4N0+huk+7+pnoXF0DsntARf9fmz1Zr1YgPIGuPWw
NxlSpG8B8on5Z7jOWQUTQOzJ4yEn+adPOAAKOtMv6vkz6goxG8XC86KMXH6TnRoj
U/5X+F2d41P8M2Qd59WZ8Q6zTp8crHFe1SF1N1oGB12ZHYDm/3lAXcgWCfOjlMDt
W7dz6iMkz8Hlun85yGQwbmzELIVp+c4jB515OEPrAYnNf2Ov9fA2VQA4aiiZERBD
d6vjnEeQXeRpJakCQ95prRmRjQkGwZbY7YQoZnmE2QyCL3THH351kjr4E+qDr8y0
McBwruo99sJ3+F4Dm1OnyDAhTNDgJNd37LRD39bxkBzCAbkVByjsMmdkAgO4s5rD
BG+Zi99JAmd6hpJR1ZPf4I7F4+sbZJYDm3hcaVNG3qbUzpw56UxM/Q/u1OMnhdAF
ICubcuyjobNWxZIHYtLXp0plUKz/CGetWwd1fv3xA9ClWN0gU5XQ5g72PcAR5Y8s
W2hZaaDJMzw62Sb38GpjarNTaLuyMk39pBNdmAynHIEWgdmvs70uBMz3hSo2HsEn
hRwKABsEI9SQZD+98rZJtXbeY5zqTeo/THT6mXl/4rs40kgwV9Hzq3/TgiiW5dvV
O2jlE7JnWDZ0S61f4yZX2MVUNSmmtHP+wEjDxMuJtGoodUP+iy7YGEZNBCm8PCM2
qjNPxoX2nearFS6dPzk23SEuHPzJRmxhtBJ7uHtaBuilBSxqRVkgRIfgYKAdHYCN
yg8o06aZZkbspOei47g6mrat/1c1tqhvEGCBfW3S+6FixdMSQr/6MAwdCst9Ud4h
l04h0peNJS9vOD7R/f1Avc0Fsgnk6BGD2RycCRjkbuz4Wnq24Yv7yFgjes2KDXi+
QflKLOaDsi0MjcRmJuJ3AYC/WlvZJb1VnQ2hgfn2bZATWV8RmBSbZB3+OvGnRM/w
KfPAh9JV1lE8+Wf1+FHXToY4V/EfI/eRz24YmhQnCrQthhohIvMFpY0g9xSjcTvv
N4Kcw5L7Z/BtZv4b4q4HonAR+ZYaFSaeeNaEY4vX0bWcK0wv4v2smqYtbrjSctX5
z6Hv6bYWAb5MGedKNvqgAJO4eP9MNx5m0b2wYm3NTNtwa+n16f+NJ36L++8TdnDh
c+DSxVxgr+VV+t+cvbJoAUM89szws5d21NNgV57rBsAB/oS6Hv8HkD70d78hbHEv
qu1Umt97T7DmRL9sDQ/i2IalV3VxsRy3seb8QS6TkqKbPI6dt5WguSS5ykJ2c7Se
svMmiIWwhODVNPiz6yStFddoC95VHnfk5BPrxY3lW664i0dtupFKBmSP756DZ4s5
uuV+d5Eb8qx/dU1J2TBEkf2HcX9B9rH490StMvmgYrOWznF8gdDoDobiA/YnXpRY
qT/7GXFDr7JcePV8yl5dyRWal0jbw+gDOfHEMHqfEbED2YWaOgs3BNg7h1IBi9wx
obaZqA8CsIU9+tvyL2PosOFGDxKoVufBDcjAPdVRWIsC65m2IKDbegxhJTI/Ab60
Fb321f0qqPQ5rnTDPGdWC8Wp0UlhCNqfRUPxZTKbJZNQSbPDXSX/8GdMzVdncjJs
jF2mThiBz3X2JXRG3FBR3CTFd8QtX5xLubt4yfZx8f/Y8wCYIZ9f48mVCXd60dZa
gJ0L2kBkO7JuQZkP5kkJfKkVsb2y6cH4Y5lH9zmILH1L86l2TLPZY/sjwpeuZwoV
V4rVsH5OHXeEXvpYvS00j7pyV9pO3aGMMwQY9d38z39ES1mFpQalJc7erDpdQpKD
i1l9MCnurgX163jkM2Xsdv3woZRAkFBYdm0Bf7J5HFe08VhEG77xHFSR9R2h0F3r
kLLfuHUaL6zxOa7+GjAj4XrQlNBEkN5cln/Vi3jOR9cdTYR0jXt+Wn+5xteSvfHz
OPhb8I08Zres7F/atSQxmTaa3l0d1sUGAt/CIbWYQxLHCPxP9YCeNT6ZngTaHoAo
NxMZO8p9Qnj6/8fMPtqR5gr3hhC9ifNNY0wugwXlvXhj1++zEUHRdPORyX0c0ebn
RqqFu6wYaPgRLixBMsVl5D6Em3MITbeKV4y2/tpL1bTcjD9aR6kYTUpg86WbtI55
UPYJV4r8Tw7HRZMmEybp+mTNfyuTCHKJJQjlJQbR2xclXPkaboRPHmatkI9r2Txk
ZqqeOX6eQ+WMO2mHW7uOFBQ5gsoiHf5PJT5XjYQmsTvashSCd+4T+7hE+Y/9x1jl
+AVGasbG/vZvGWF6GoWgxTNkOOTx+1q8fyUTC/aolK2v1h7nFKHqx9Oht+15EFJL
FciCcaNJ7i46Uwq3+lUnoan22doRtmbIcRqYLCzL0dHlEPQaaUgNSeCeXYMttZt5
o+o/96QxkfQdDDmBVNIQF6XdKXUBqtgEnUu3jadKVnnj6rV7tN2xSUz1HoGKnpVJ
oaCvL148MB8XT7JSW5gXOVqSt0ygrYttzLG+u+TliLwTHUED4SfQ6O52J/6jXnd6
kbykHvfbyn3PadTlg82A4H18kztYzkq3WSyKM9Y6SmJrdb+Im+9/GbIuc5v1VMez
b1fay1S2NFs2xyg52fkm6P+/IcTY9ji+XHQLf6uC1GSSI+KehIrqd/93yU3phT3P
aQqRLKEBo8cAorugqD9c/poooUF9tBc9iqqkH9NK45EocCQRSbyqq8ewBR2H/yOu
R0hF/+AKHCnZG8iLQXCrBBfYsy4tncQorH8C3w2SGWCCJDUt7im/Chqk8A2XG+Y5
XP0K6G2G/YbNugOGBOTt38TMi6Hyv/SoBQSln0+uqc3DinOXcH7qQDV1pkM0mSoH
80KDJDwojFX6WEEw+LcBijf1B0s051TbwII9561f+WYEA2odKuOSpKm/rt36nvSh
SDpkj2uvnmb7RnpCYsw+cXn9ZxTv36eVuOwub/8iWoRDGGfRuKaQvcG0MraYjn0V
hYNxQQxnkfnFqPNR7e6Cw1wSRJXnFw0zntoVmYBcp+H0bNmzWM2DCbb++pThxZrS
9TeL1q2OAZAKhMJunxQ/eiIOX7KBMut70PhMMVMasH7O583h/LjApdtXe43qdX3g
iesoR7OVavput3UE3QUBKykByUIOYHzFRlp2sOHFvlldivhBJ60KY0BUQxDlHzaa
CLGvgMPdJ3vahmbTfxyQZx1bco/AmaL02PM1Cw7ZfVvuWtdwyst+qSlLJ68ZVCN6
2YFTZmn0DkVcZgEeOyMpThYZAeWdR8Gd5VfFVB4jzG2VbudC23CgKAg0MroY70zX
JwF+oIYtnkW5d6ip27ANXemD6wJDrZIlE0ZW2kv/rZeN6e9wuzskhZekJanMZMHb
WSj+nIzIpbyi7dCtu+uEB3OIEAehXOVT2vV8nHFia1U1J9jYUduUfIVc7MGS3I+f
tVVzdcz3OvZtUFRzsbbRZNOkTYbdDldIg00Dqsx614qNiBlA9QO9MBXlfTK9XzeZ
EVr71euMZ2OVK5dg69+n0Pr2KknuldnQNIqTedLrv7lnLYHZYcrOtBuh+Q63iNEb
ZRwQb63weIDTNkeqIfLRFWLBIBVKjCoZufWDJA+4Aa8FTJbOlcZlIEP2ukke7uUg
67wykpKEB1emqy1kFjRGzbhp9yWrf5cxKB81dGh12gDhg4r7eHTAVh+zbKugwsVy
r2+6ew/8rV5rolw4vpIsf9omPEZQyVtIYZOCXOBFUdr0fkTFdJdmd+tLW+EZG2A0
NrwXItt9Kr4NJoQCkFhd+CJ7rUVDYSNrFPDS43k0JVQnjoH5NHS+bRhdlv0ieQNH
ZygmYarLM5/aGoSw7mbtBJ2FK4Yu51HOeb+YpM2EpaGOfc0f1yATDbXFLvNmr42C
5hOip+gF9cjQ8yar91y+x7L4cScJlAP/15N36ZOQvUon5U7/Q2YH6zgm5STeorkT
A2sHqBnDzzolnbPjwDfB9YrIeImkRUbOID22+aUAQm+BBhwGJfQsHWZk/QC4wj5U
9FVU6Gso41QUnusQmJ5uxBXJ8X9DewNsXXGQZCvgg4EF3y4S6UtcaFew6u6iXKIk
ggGpSBiFSQodOHlXhpck2ppmDidBuxLimCscEiqsn1JzC2UQjdNdgsa2SmOZ5vt7
8tNfeQ4rhhBcipj25rneji3k9+E9YzwDy7ow4x3hNUCSzm+unZn6aIyOgzLCGI48
6/xT/e97sWRBpTYehnsbhSVLKZle/Fmno8qrLtbVNIT2v3sw/n1OMa1i63VXS2L0
eplX1T76hiIvT+gF6wskN2Y8YafocCRaf0XNBRjb69aRRdy2vAtIwUHqjjz1k0Ez
lts24SVV0o4fjMj/7c4qJzJIdd4Aqw/1g8xYLL8Mu7An3hpjfOR1uzH/5WZIGjbC
5Z4RZuzGoHD2xmwkl8putm5h4XV74uaFz5n3vsgSOd59+dWUw0hkjD8KtDoml7sd
Gsu3DMwgq0iu2sLLyuwPgTvfYPwKRmQSGQl/fL6qMCCXeAEh+u++amyYSvPlXsm6
SryPZHwBF2fRXzN33cOo3RWYPIsHMtHkz4le2WgOLjpxm82SAp5+DP0hXZf+j2O+
Gf5oZwzBhqXnRG66T8FZ5LX2DHXM9245FiJ42IuXP+WwSLQVmjM6BDeZegAmj5WA
zfpeMDB87bhgAIpLHWjf/VOWS9FTDMq5j2oM76VGVnvYvHo+Tjt9TMFFXAvNGEuJ
WKfhEgb7lobBV8Fwej2gD8N1gAY+7tOSLDcAycNTCX0AI/Hpyf10ykirGQcuAmiK
zNZdcT9Oj07vgO5vqNglw8fEO4Tnd7ngqg45sXX7eo73fKoFR7X7adxuAHPdjwPl
DI06RjSv1z+TbuxQZw0eISBslc8OX3GRoLGM2amPeHwNFXlg9jQdW7DSmIxlTTug
XhplEe0d1CNHie3t2MxkU5NpygUDkEV0jfcVkGBrYFVTsbyHNepdwCH1x248QiTm
NtvuRtJki3lO1iFsx9D8duoBlBKpoE+0mNalcB+nywFH2ujfiRptB3wr7zQT7GwB
RDpgT0+aGoZGL2m9LMYsgfKev039C0nMEBT4p0uw1c1QFtva5p1amvVgG9X/4cEz
Y+25I1qEcGE4lq+xMHG5eSG+XjDOhDvrq6K0NTrhq5EaDyjAuZRV/R0MfApb7JQq
dTwBFRc/uHnW1xi/wofYL+U9bvAg9s6oeiz70VVewOzEBXIQDiYhH4rys9xLhRih
ccyg796PR+LWWjIHKMLjFTptWxVEoP1RxPTn/Sg4B9Vys+lVkT/ua+AtjbSfPPnc
C4m09/EO6CPiIqIlMw8CySCcoXuzj/KIxbvdzRD4M0dXAkc/dAjU2/kJGtb6chTV
iMZvELImu9pTp9na+AVcQvuc7yChd44+YrIeZLTPTf4Pr+2UwgMrfZuZK5CWhmDb
+x/aLvVWVDLnCLZBp06eGqbdREEziiCglki5B08C0XsHwXC/s5/mx1j13OedWZUO
2btQxDfhB0IAS8RWRdp8u1LQEC5PM3G7uHE1/wDuhs4E7x4d4ea4K4Wmk7xd02Sv
Z96zdlfzGjDxUj2hY4N0F4kI4VAQaanClKaSHJaODsO93GYDbim0jvWdx5Ed8A8F
HmMRk4ocGjzA+7nLu70eEpXZfyc2Ch/xXAbUvIr2M7aXluPJ0mcyCjr5HakxWBF9
A8fP5T+4MZZ78y5lqkagDmvQFCBY3RW8Qsfw0TjQsGeUYh6GqkXkU9PSxge/CWHN
bY71ZkTgPJK3g5Re9nynjBi1+N0BHriMuOG7s2L5Ao6JNp2eXTm1wTBUXpdvZy9g
+E/ET8x9nQ8o3eQLs5o6x6wFCr5btDiOgJn/2J7crBZL6hFAG75CLLKxM5n6qSei
hE7LDLuAK3hLW3XyYAh0wnt1j64WqTjiSyv5+FVgEjUaA+QBy+w+ytKDLbjgXen/
Vn3fmqeNnCdH/+vMMcYoItxyF0qDEpaan+obuJOr5/0Hq5eZDeZ+jRDaRS9B9tsz
QmsJYDsnr4DALN2BZfLl89OoLXOOfPeaA7mtUi2g/3cAxDPCTHNXAGxwIqUnOWvJ
bIcHIqWszg4be/zRIzgV2mCVKmh4vXCpS0mFFdIsjY2cW5SG77cAjVySns66kCZE
nWuAvENiEeuE08uUq+Y3qq413KFH5IRhcTdrkxpONT6eg4QbNq7cS1ERoYcPORLl
t8cVGF8/B6U0E2H0IMQ4nBE4962SfE5quXMxj4IBM0goEUkhKptn99HSzkUxobcM
sJ2vTVyrjw5+Jc4Wl90L4VHjU0Wb1AzMMk9t/T7e0KOs7BpjsO2g0gKNssgYVnxM
CJknn7VsVnhvAL1nf14JCw==
`pragma protect end_protected