/*******************************MILIANKE*******************************
*Company : MiLianKe Electronic Technology Co., Ltd.
*WebSite:https://www.milianke.com
*TechWeb:https://www.uisrc.com
*tmall-shop:https://milianke.tmall.com
*jd-shop:https://milianke.jd.com
*taobao-shop1: https://milianke.taobao.com
*Create Date: 2019/12/17
*Module Name:
*File Name:
*Description: 
*The reference demo provided by Milianke is only used for learning. 
*We cannot ensure that the demo itself is free of bugs, so users 
*should be responsible for the technical problems and consequences
*caused by the use of their own products.
*Copyright: Copyright (c) MiLianKe
*All rights reserved.
*Revision: 1.0
*Signal description
*1) I_ input
*2) O_ output
*3) IO_ input output
*4) _n activ low
*5) _dg debug signal 
*6) _r delay or register
*7) _s state mechine
*********************************************************************/
`timescale 1ns / 1ns

/*uiphyrst ��λ�������*/

module uiphyrst#
(
parameter integer  CLK_FREQ = 32'd100_000_000         //ʱ�Ӳ���
)                                            //���÷�Ƶϵ����������ˮ�Ƶı仯�ٶ�
(                                            //�ò����������ϲ����ʱ�޸�
 input   wire       I_CLK,                   //ϵͳʱ���ź�
 input   wire       I_rstn,                  //ȫ�ָ�λ
 input   wire       I_phyrst,                //��λʱ��
 output  reg        O_phyrst,                 //��λ���
 output  wire       O_phyrst_done
);

localparam  T_SET = CLK_FREQ/100;

reg [31:0] t_cnt; //100ms ������
reg [1 :0] S_PHYRST;

reg  phyrst_r1,phyrst_r2,phyrst_r3;
reg  phy_rst_req; //��λ����
wire phy_rst_done = (S_PHYRST == 3);//��λ���
wire phy_rst_ack  = (t_cnt == T_SET);//��λ������Ӧ��

assign O_phyrst_done =   ~phy_rst_req&I_rstn;      

always @(posedge I_CLK )begin //ץȡ��λ
    phyrst_r1  <= I_phyrst;
    phyrst_r2  <= phyrst_r1;
    phyrst_r3  <= phyrst_r2;
end

always @(posedge I_CLK or negedge I_rstn)begin
    if((I_rstn == 1'b0) || ({phyrst_r3,phyrst_r2} == 2'b01)) //�ϵ縴λ���ߴ�����λ
       phy_rst_req <= 1; 
    else if(phy_rst_done)   //ϵͳ��λ,����PHY��λ���
       phy_rst_req <= 0;    
end

//PHY��λ��������󣬼���������
always @(posedge I_CLK)begin                                       
    t_cnt <= phy_rst_req ?  
             phy_rst_ack ? 0 : t_cnt + 1'b1
             : 0 ;  
end

//��λ״̬��
always @(posedge I_CLK or negedge I_rstn)begin
    if(I_rstn == 1'b0 )                             
       S_PHYRST <= 0;   
    else begin
        case(S_PHYRST)
        0:if(phy_rst_req) S_PHYRST <= 1;//��λ��ʼ
        1:if(phy_rst_ack) S_PHYRST <= 2;//�͵�ƽ20MS
        2:if(phy_rst_ack) S_PHYRST <= 3;//�ߵ�ƽ20MS
        3:S_PHYRST <= 0;//��λ���
        default :S_PHYRST <= 0;
        endcase
    end
end

//����100MS ���帴λ
always @(posedge I_CLK)begin
    if(S_PHYRST == 2) O_phyrst <= 0;
    else O_phyrst <= 1;
end

endmodule   

