

`timescale 1ns / 1ns

module uicfg_imx415#
(
parameter	 CLK_DIV  = 16'd999
)
(
input  wire             I_clk,  //ϵͳʱ������
input  wire             I_rst_n,  //ϵͳ��λ����
input  wire             I_ae_req,//����ͷAE����
input  wire	 [7:0] 		I_ae_data,
output wire             O_cam_scl, //I2C���ߣ�SCLʱ��
inout  wire             IO_cam_sda, //I2C���ߣ�SDA����
output reg              O_cfg_done, //�������
output reg              O_ae_cfg_done
);	

localparam CAM_ID = 8'h34;//������ַ 

reg  [7:0] rst_cnt;//��λ��ʱ����
reg  [21:0] cnt;//����ģʽ�Ĵ�����ʱ���ü���

reg  O_cfg_done_r;//����ģʽ�Ĵ�����������ź�
reg  iic_req;//�������I2C�������ź�
wire ic_busy; //I2C������æ�ź� 
wire   O_iic_bus_error;
reg  [31:0] wr_data;     //д���ݼĴ���
reg  [1 :0] TS_S = 2'd0; //״̬���Ĵ���
reg  [7 :0] reg_index;   //�Ĵ�����            
                                             
reg [23:0] REG_DATA;    //�Ĵ�������
reg [7:0]  REG_SIZE;    //�Ĵ�������

wire [23:0] REG_DATA_REG; //�Ĵ�������
reg  [23:0] REG_DATA_ST;  //�����Ĵ�������
reg  [23:0] REG_DATA_AE;  //AE�Ĵ�������

wire [7 :0] REG_SIZE_REG; //�Ĵ�������
wire [1 :0] REG_SIZE_ST = 2'd2;  //�����Ĵ�������
wire [2 :0] REG_SIZE_AE = 3'd4;  //AE�Ĵ�������


//�ڲ�����������һ���ӳٸ�λ
always@(posedge I_clk or negedge I_rst_n)  
    if(I_rst_n == 1'b0) //��λ��ʼ���Ĵ���
        rst_cnt<= 8'd0; 
    else if(rst_cnt[7] == 1'b0)
       rst_cnt <= rst_cnt + 1'b1; 
    else 
       rst_cnt <= rst_cnt; 
	   
always@(posedge I_clk or negedge I_rst_n)  begin
    if(I_rst_n == 1'b0) //��λ��ʼ���Ĵ���
         cnt <= 0;
    else if(cnt == 1000_000)
         cnt <= 0;
    else if(O_cfg_done == 1'b1)
         cnt <= cnt + 1;
    else if(O_cfg_done_r == 1'b1)
         cnt <= cnt;
end

always@(posedge I_clk or negedge I_rst_n)begin
    if(I_rst_n == 1'b0)begin
		REG_SIZE <= 8'b0;
		REG_DATA <= 24'b0;
	end
	else if(O_cfg_done == 1'b0)begin
		REG_SIZE <= REG_SIZE_REG;
		REG_DATA <= REG_DATA_REG;
	end
	else if(O_cfg_done == 1'b1 && O_cfg_done_r == 1'b0)begin
		REG_SIZE <= REG_SIZE_ST;
		REG_DATA <= REG_DATA_ST;
	end
	else if(O_cfg_done == 1'b1 && O_cfg_done_r == 1'b1)begin
		REG_SIZE <= REG_SIZE_AE;
		REG_DATA <= REG_DATA_AE;
	end
	else begin
		REG_SIZE <= 8'b0;
		REG_DATA <= 24'b0;
	end
end

always@(posedge I_clk ) begin 
    if(rst_cnt[7] == 1'b0)begin //��λ��ʼ���Ĵ���
        reg_index  <= 9'd0;
        iic_req    <= 1'b0;
        wr_data    <= 32'd0;
        O_cfg_done <= 1'b0;
        O_cfg_done_r <= 1'b0;
        O_ae_cfg_done <= 1'b1;
        TS_S     <= 2'd0;    
    end
    else begin
        case(TS_S)
        0:if(reg_index == REG_SIZE && O_cfg_done == 1'b0) begin//����������
            O_cfg_done <= 1'b1;       //���� cfg_done��׼
        end 
        else if(reg_index == REG_SIZE && O_cfg_done == 1'b1 && O_cfg_done_r == 1'b0) begin//����������
            O_cfg_done_r <= 1'b1;       //���� cfg_done��׼
        end 
        else if(cnt== 1000_000)begin
            O_cfg_done_r <= 0;
            reg_index   <= 0;
        end
		else if(reg_index == REG_SIZE && O_cfg_done == 1'b1 && O_cfg_done_r == 1'b1) begin//����������
            O_ae_cfg_done <= 1'b1;       //���� cfg_done��׼
        end 
        else if(I_ae_req)begin
            O_ae_cfg_done <= 0;
            reg_index   <= 0;
        end
        else if((O_cfg_done&O_cfg_done_r&O_ae_cfg_done) == 1'b0)
            TS_S <= 2'd1;           //��һ��״̬
        1:if(!iic_busy)begin        //�����߷�æ���ſ��Բ���I2C������
            iic_req  <= 1'b1;       //�������I2C������
			wr_data[7  :0] <= CAM_ID;           //������ַ   
			wr_data[15 :8] <= REG_DATA[23:16];  //�Ĵ�����ַ-��8bit    
			wr_data[23:16] <= REG_DATA[15: 8];  //�Ĵ�����ַ-��8bit  
            wr_data[31:24] <= REG_DATA[7 : 0];  //�Ĵ�������
            TS_S      <= 2'd2; //��һ��״̬
        end    
        2:if(iic_busy)begin
             iic_req  <= 1'b0;  //���� iic_req =0
             TS_S     <= 2'd3;  //��һ��״̬
        end
        3:if(!iic_busy)begin  //�����߷�æ���ſ��Բ���I2C������ 
			reg_index<= reg_index + 1'b1;//�Ĵ���������1
			TS_S    <= 2'd0;//�ص���ʼ״̬
        end 
        endcase
   end
end

//����I2C����ģ��
uii2c#
(
.WMEN_LEN(4),     //���֧��һ��д��4BYTE(����������ַ)
.RMEN_LEN(1),     //���֧��һ�ζ���1BYTE
.CLK_DIV(CLK_DIV) //100KHZ I2C����ʱ��
)
uii2c_inst
(
.I_clk(I_clk),//ϵͳʱ��
.I_rstn(rst_cnt[7]),//ϵͳ��λ
.O_iic_scl(O_cam_scl),//I2C SCL����ʱ��
.IO_iic_sda(IO_cam_sda),//I2C SDA��������
.I_wr_data(wr_data),//д���ݼĴ���
.I_wr_cnt(8'd4),    //��Ҫд������BYTES
.O_rd_data(),       //�����ݼĴ���
.I_rd_cnt(8'd0),    //��Ҫ��������BYTES
.I_iic_mode(1'b0),  //��ģʽ����
.I_iic_req(iic_req),//I2C����������
.O_iic_busy(iic_busy),//I2C������æ
.O_iic_bus_error(O_iic_bus_error)
);


//����CAM�ļĴ������ñ�
uiimx415reg uiimx415reg_inst
(
.REG_SIZE(REG_SIZE_REG),  //�Ĵ�������
.REG_INDEX(reg_index),    //�Ĵ�����
.REG_DATA(REG_DATA_REG)   //�Ĵ�������
);  

always@(*)
   case(reg_index)
		0:		REG_DATA_ST = {16'h3000, 8'h00}; 
		1:		REG_DATA_ST = {16'h3002, 8'h00}; 
		default:REG_DATA_ST = {16'h0000, 8'h00};
   endcase

always@(*)
   case(reg_index)
		0:		REG_DATA_AE = {16'h3090, I_ae_data}; 
		1:		REG_DATA_AE = {16'h3092, I_ae_data}; 
		2:		REG_DATA_AE = {16'h3094, I_ae_data}; 
		3:		REG_DATA_AE = {16'h3096, I_ae_data}; 
		default:REG_DATA_AE = {16'h0000, 8'h00};
   endcase

endmodule
