module cwc5
(
  input   [0:0]                 probe0,
  input   [0:0]                 probe1,
  input   [0:0]                 probe2,
  input   [8:0]                 probe3,
  input   [8:0]                 probe4,
  input   [15:0]                probe5,
  input   [0:0]                 probe6,
  input   [15:0]                probe7,
  input   [0:0]                 probe8,
  input   [0:0]                 probe9,
  input   [0:0]                 probe10,
  input   [0:0]                 probe11,
  input   [15:0]                probe12,
  input   [0:0]                 probe13,
  input   [0:0]                 probe14,
  input   [7:0]                 probe15,
  input   [8:0]                 probe16,
  input   [15:0]                probe17,
  input   [15:0]                probe18,
  input   [0:0]                 probe19,
  input   [0:0]                 probe20,
  input   [0:0]                 probe21,
  input   [3:0]                 probe22,
  input   [15:0]                probe23,
  input   [0:0]                 probe24,
  input   [3:0]                 probe25,
  input   [0:0]                 probe26,
  input   [8:0]                 probe27,
  input   [15:0]                probe28,
  input   [30:0]                probe29,
  input   [0:0]                 probe30,
  input   [15:0]                probe31,
  input   [0:0]                 probe32,
  input   [255:0]               probe33,
  input   [0:0]                 probe34,
  input   [0:0]                 probe35,
  input   [30:0]                probe36,
  input   [0:0]                 probe37,
  input   [15:0]                probe38,
  input   [0:0]                 probe39,
  input   [255:0]               probe40,
  input   [0:0]                 probe41,
  input   [0:0]                 probe42,
  input                         clk
);

  ChipWatcher_04b294874e40  ChipWatcher_04b294874e40_Inst
  (
      .probe0(probe0),
      .probe1(probe1),
      .probe2(probe2),
      .probe3(probe3),
      .probe4(probe4),
      .probe5(probe5),
      .probe6(probe6),
      .probe7(probe7),
      .probe8(probe8),
      .probe9(probe9),
      .probe10(probe10),
      .probe11(probe11),
      .probe12(probe12),
      .probe13(probe13),
      .probe14(probe14),
      .probe15(probe15),
      .probe16(probe16),
      .probe17(probe17),
      .probe18(probe18),
      .probe19(probe19),
      .probe20(probe20),
      .probe21(probe21),
      .probe22(probe22),
      .probe23(probe23),
      .probe24(probe24),
      .probe25(probe25),
      .probe26(probe26),
      .probe27(probe27),
      .probe28(probe28),
      .probe29(probe29),
      .probe30(probe30),
      .probe31(probe31),
      .probe32(probe32),
      .probe33(probe33),
      .probe34(probe34),
      .probe35(probe35),
      .probe36(probe36),
      .probe37(probe37),
      .probe38(probe38),
      .probe39(probe39),
      .probe40(probe40),
      .probe41(probe41),
      .probe42(probe42),
      .clk(clk)
  );
endmodule
