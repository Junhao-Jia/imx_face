
/*******************************MILIANKE*******************************
*Company : MiLianKe Electronic Technology Co., Ltd.
*WebSite:https://www.milianke.com
*TechWeb:https://www.uisrc.com
*tmall-shop:https://milianke.tmall.com
*jd-shop:https://milianke.jd.com
*taobao-shop1: https://milianke.taobao.com
*Create Date: 2023/08/07
*Module Name:key
*File Name:key.v
*Description: 
*The reference demo provided by Milianke is only used for learning. 
*We cannot ensure that the demo itself is free of bugs, so users 
*should be responsible for the technical problems and consequences
*caused by the use of their own products.
*Copyright: Copyright (c) MiLianKe
*All rights reserved.
*Revision: 1.0
*Signal description
*1) I_ input
*2) O_ output
*3) IO_ input output
*4) S_ system internal signal
*5) _n activ low
*6) _dg debug signal 
*7) _r delay or register
*8) _s state mechine
*********************************************************************/
`timescale 1ns / 1ns
module key #
(
parameter REF_CLK = 64'd50_000_000        //����ʱ��Ϊ�����������ϲ�����޸�
)
(
input  I_sysclk,
input  I_rstn,
input  I_key,
output O_key_down,
output O_key_up
);

parameter  T10MS = (REF_CLK/100 - 1'b1);                      //����10MS��ʱ�ӷ�Ƶ����
parameter  KEY_S0 = 2'd0;                                      //���ð���״̬����״̬
parameter  KEY_S1 = 2'd1;
parameter  KEY_S2 = 2'd2;
parameter  KEY_S3 = 2'd3;

reg [32:0] t10ms_cnt = 25'd0;
reg [3:0] key_r = 4'd0;
reg [1:0] key_s = 2'b0;
reg [1:0] key_s_r = 2'b0;
wire t10ms_done ;
 
assign t10ms_done = (t10ms_cnt == T10MS);
assign O_key_down   = (key_s == KEY_S2)&&( key_s_r == KEY_S1);    //�����жϰ�������ʱ������
assign O_key_up     = (key_s == KEY_S0)&&( key_s_r == KEY_S3);     //�����жϰ����ɿ�ʱ������

//10ms timer counter
always @(posedge I_sysclk or negedge I_rstn)begin                 //ϵͳʱ�ӵ��������Լ���λ���½��ش���
    if(I_rstn == 1'b0)begin
        t10ms_cnt <= 25'd0;                                          //ϵͳ��λ
    end
    else if(t10ms_cnt < T10MS)                                        //10ms������Ŀ��ֵ�� T10MS
        t10ms_cnt <= t10ms_cnt + 1'b1;                                //δ�ﵽĿ��t10ms_cnt+1 
    else 
        t10ms_cnt <= 25'd0;                                             //�ﵽĿ��ֵ��λ
end
always @(posedge I_sysclk)begin                                     //��key_s��״̬����һ��
    key_s_r <= key_s;
end
always @(posedge I_sysclk)begin                                     //��I_key��״̬����һ��
    key_r <= {key_r[2:0],I_key};
end
always @(posedge I_sysclk or negedge I_rstn)begin                //����״̬�����趨������4��״̬
    if(I_rstn == 1'b0)begin
        key_s <= KEY_S0;
    end
    else if(t10ms_done)begin                                           //��������Ϊt10ms_done��˵���������е�״̬ת�ƶ���ÿ10ms
        case(key_s)                                                     //����һ��
            KEY_S0:begin
            if(!key_r[3])                                                //�յ���һ�������ĵ͵�ƽ�źţ������ж��Ƿ�Ϊë��
                key_s <= KEY_S1;                                        //ת��״̬S1
            end  
            KEY_S1:begin//recheck key done                               //�ڶ����жϰ����Ƿ���
            if(!key_r[3])
                key_s <= KEY_S2;                                        //����ת��S2״̬
                else 
                key_s <= KEY_S0;                                        //û���£��ж�Ϊë�̣�ת��S0״̬���ȴ�����
            end 
            KEY_S2:begin//wait key up                                     //ȷ���������º�
            if(key_r[3])                                                //�ȴ������ɿ������յ������ĸߵ�ƽ�źţ�
                key_s <= KEY_S3;                                        //����ȷ���Ƿ�Ϊë��
            end                                                              //ת��״̬S3
            KEY_S3:begin//recheck key up                                   
            if(key_r[3])                                                 //�ڶ����жϰ����Ƿ��ɿ�
                key_s <= KEY_S0;                                           //��Ȼ��⵽�������ɿ���״̬��ת��S0״̬���ȴ�����
            end
        endcase                  
    end
end

endmodule   
