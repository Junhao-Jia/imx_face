/*****************************************************************
Company : MiLianKe Electronic Technology Co., Ltd.
WebSite:https://www.milianke.com
TechWeb:https://www.uisrc.com
tmall-shop:https://milianke.tmall.com
jd-shop:https://milianke.jd.com
taobao-shop: https://milianke.taobao.com
Description: 
The reference demo provided by Milianke is only used for learning. 
We cannot ensure that the demo itself is free of bugs, so users 
should be responsible for the technical problems and consequences
caused by the use of their own products.
@Author      :   XiaoQingquan 
@Time        :   2024/10 
version:     :   
@Description :   ��ԭ������ɾȥ��һЩ׸��Ĵ��룬�����Ż���ʱ�򣬼���BRAM IP�ˣ�
                 �ôӳ�����������ÿһ�����ݶ����Զ�����Ӧ���������ݽ������棬ʹ
                 �����������и��ӹ㷺�ˡ�
*****************************************************************/
module awb  #(   
    parameter IMG_HEIGHT = 1080,
    parameter IMG_WIDTH  = 1920
) 
(
    input                   I_clk  ,
    input                   I_rst_n,


    input                   I_tlast  ,
    input                   I_tuser  ,
    input [95:0]            I_tdata  ,
    input                   I_tvalid , 
    output                  I_tready ,

    output                  O_tlast  ,
    output                  O_tuser  ,
    output [95:0]           O_tdata  ,
    output                  O_tvalid ,
    input                   O_tready
);


/*****************************************************************
                          �м��ź�                                        
*****************************************************************/

reg         I_tvalid_r0,I_tvalid_r1;          // ������Ч�źŵļĴ�
reg  [95:0] I_tdata_d0,I_tdata_d1,I_tdata_d2; // �������ݵļĴ�

// �ۼ�RGBͨ������ֵ�����ڼ���ƽ��ֵ
reg  [31:0]         sum_r;
reg  [31:0]         sum_g;
reg  [31:0]         sum_b;

wire  [95:0]        data_d0 ;     // ��ʱ�������
wire                valid_d0;     // ��ʱ�����Ч�ź�
wire                I_tuser_r0;   // ��ʱ���֡��ʼ�ź�

reg                 I_tuser_r1;   // ֡��ʼ�źŵļĴ�

reg   [95:0]        data_d1 ;     // �ٴ���ʱ�������
reg                 valid_d1;     // �ٴ���ʱ�����Ч�ź�
reg   [9:0]         rgb_sum;//ÿ�����ص�RGB�ĺ�
localparam IMG_WIDTH_4x = (IMG_WIDTH >> 2);  // ͼ���ȳ���4���õ�ÿ�����ݿ������

/*****************************************************************
                           ƽ��ֵ����                                        
*****************************************************************/

// ���������ݺ���Ч�źŽ��мĴ棬�γ���ˮ��
always @(posedge I_clk or negedge I_rst_n) begin
    if (!I_rst_n) begin
        I_tdata_d0  <= 0;
        I_tdata_d1  <= 0;
        I_tdata_d2  <= 0;
        {I_tvalid_r0,I_tvalid_r1} <= 0;
    end else begin
        I_tdata_d0  <= I_tdata   ;
        I_tdata_d1  <= I_tdata_d0;
        I_tdata_d2  <= I_tdata_d1;
        I_tvalid_r0 <= I_tvalid;
        I_tvalid_r1 <= I_tvalid_r0;
    end
end


// ���������ݲ��Ϊ4�����ص�RGB����
wire [7:0] rgb888_r_d;
wire [7:0] rgb888_g_d;
wire [7:0] rgb888_b_d;

assign  rgb888_r_d = I_tdata[16+:8];
assign  rgb888_g_d = I_tdata[8+:8];
assign  rgb888_b_d = I_tdata[0+:8];


// ���������ݲ��Ϊ4�����ص�RGB����
wire [7:0] rgb888_r_d0;
wire [7:0] rgb888_g_d0;
wire [7:0] rgb888_b_d0;

assign  rgb888_r_d0 = I_tdata_d0[16+:8];
assign  rgb888_g_d0 = I_tdata_d0[8+:8];
assign  rgb888_b_d0 = I_tdata_d0[0+:8];


    ///������ɫ
    always @(posedge I_clk or negedge I_rst_n) begin
        if(!I_rst_n) begin
            rgb_sum <= 0;
        end
        else if(I_tvalid)begin
            rgb_sum <= rgb888_r_d + rgb888_g_d + rgb888_b_d;
        end
    end
    
    wire flag_frame_r;
    reg [31:0] sum_r_d ;
    reg [31:0] sum_g_d ;
    reg [31:0] sum_b_d ;
    // ��ÿ��ͨ����ֵ�����ۼӣ����ڼ���ƽ��ֵ
    always @(posedge I_clk or negedge I_rst_n) begin
        if (!I_rst_n ) begin
            // ��λ���п�ʼ�ź���Чʱ�������ۼ���
            sum_r <= 1;
            sum_g <= 1;
            sum_b <= 1;
        end else if (flag_frame_r) begin
            // ��������Чʱ���ۼ�RGB������ֵ
            sum_r <= sum_r_d;
            sum_g <= sum_g_d;
            sum_b <= sum_b_d;
        end else if (I_tvalid_r0 && (rgb_sum < 700)) begin
            // ��������Чʱ���ۼ�RGB������ֵ
            sum_r <= sum_r + rgb888_r_d0;
            sum_g <= sum_g + rgb888_g_d0;
            sum_b <= sum_b + rgb888_b_d0;
        end
    end

    reg [3:0]  frame_cnt;
    always @(posedge I_clk or negedge I_rst_n) begin
        if (!I_rst_n ) begin
            sum_r_d <= 1;
            sum_g_d <= 1;
            sum_b_d <= 1;
        end else if(frame_cnt==4)begin
            sum_r_d <= 1;
            sum_g_d <= 1;
            sum_b_d <= 1;
        end else if(I_tvalid_r0 && (rgb_sum < 700))begin
            sum_r_d <= sum_r_d + rgb888_r_d0;
            sum_g_d <= sum_g_d + rgb888_g_d0;
            sum_b_d <= sum_b_d + rgb888_b_d0;
        end 
    end

    always @(posedge I_clk or negedge I_rst_n) begin
        if (!I_rst_n ) begin
            frame_cnt <= 0;
        end else if(frame_cnt==4)begin
            frame_cnt <= 0;
        end else if(I_tuser)begin
            frame_cnt <= frame_cnt + 1;
        end
    end

    reg  flag_frame;
    always @(posedge I_clk or negedge I_rst_n) begin
        if (!I_rst_n ) begin
            flag_frame <= 0;
        end else if(frame_cnt==1)begin
            flag_frame <= 1;
        end else begin
            flag_frame <= 0;
        end
    end


    reg  flag_frame_d;
    always @(posedge I_clk or negedge I_rst_n) begin
        if (!I_rst_n ) begin
            flag_frame_d <= 0;
        end else begin
            flag_frame_d <= flag_frame;
        end
    end

    assign flag_frame_r = (flag_frame == 1) && (flag_frame_d == 0);



  /*****************************************************************
                           ��������                                       
*****************************************************************/

  wire [47:0] dout_R;
  wire [47:0] dout_B;

  wire done;

  wire [47:0] in_r_x1;
  wire [47:0] in_b_x1;
  assign in_r_x1 = dout_R[47:0];
  assign in_b_x1 = dout_B[47:0];

    

/*****************************************************************
                   IP ����                                    
*****************************************************************/
    //Ϊ�˱�֤������ӳ٣�����ʹ���˳�����


      divider div_gen_G_R_r1 (
          .clk(I_clk),  // input wire aclk
          .rst(!I_rst_n),
          .start(I_tvalid_r1),
          .denominator(sum_r),  // input wire [31 : 0] s_axis_divisor_tdata
          .numerator({sum_g,16'd0}),  // input wire [47 : 0] s_axis_dividend_tdata
          .quotient(dout_R),  // output wire [79 : 0] m_axis_dout_tdata
          .done(done)
      );

      divider divide_G_B_r1 (
          .clk(I_clk),  // input wire aclk
          .rst(!I_rst_n),
          .start(I_tvalid_r1),
          .denominator(sum_b),  // input wire [31 : 0] s_axis_divisor_tdata
          .numerator({sum_g,16'd0}),  // input wire [47 : 0] s_axis_dividend_tdata
          .quotient(dout_B),  // output wire [79 : 0] m_axis_dout_tdata
          .done()
      );

     
    signal_delay #(
        .IMG_HEIGHT   (IMG_HEIGHT),
        .IMG_WIDTH    (IMG_WIDTH ),
        .DATA_WIDTH   (96  ),
        .DELAY_CYCLE  (50)
    )signal_delay_d (
        /*input                       */ .I_clk  (I_clk  ),
        /*input                       */ .I_rst_n(I_rst_n),
        /*input                       */ .I_tuser(I_tuser),  //synthesis keep 
        /*input  wire                 */ .I_valid(I_tvalid_r1),  //synthesis keep 
        /*input  wire [DATA_WIDTH-1:0]*/ .I_data (I_tdata_d1 ),   //synthesis keep 
        /*output wire                 */ .O_valid(valid_d0   ),  //synthesis keep 
        /*output wire [DATA_WIDTH-1:0]*/ .O_data (data_d0    ),   //synthesis keep 
        /*output wire                 */ .O_tuser(I_tuser_r0 )
    );

    

/*****************************************************************
                            ????????                                      
*****************************************************************/

reg  [19:0]   in_r_r1;
reg  [19:0]   in_b_r1;


// �������棬��ֹ������������������0xFFFFF
always @(posedge I_clk or negedge I_rst_n)begin 
    if(!I_rst_n || I_tuser)begin
        in_r_r1 <= 20'h10000;
        in_b_r1 <= 20'h10000;
    end
    else if(done)begin
        if(|in_r_x1[47:20])        // �жϸ�λ�Ƿ���1����ֹ���
            in_r_r1 <= 20'hfffff;
        else 
            in_r_r1 <= in_r_x1[19:0];
        if(|in_b_x1[47:20])
            in_b_r1 <= 20'hfffff;
        else 
            in_b_r1 <= in_b_x1[19:0];
    end
end
    ////�ź�ͬ��
    always @(posedge I_clk or negedge I_rst_n) begin
      if (!I_rst_n) begin
          valid_d1 <= 0;
          data_d1  <= 0;
          I_tuser_r1 <= 0;
      end else begin
          valid_d1 <= valid_d0;
          data_d1  <= data_d0 ;
          I_tuser_r1 <= I_tuser_r0;
      end
    end
/*****************************************************************
                           ????????                                       
*****************************************************************/

    reg [27:0] R_new_r1;
    reg [27:0] G_new_r1;
    reg [27:0] B_new_r1;

    reg [27:0] R_new_r2;
    reg [27:0] G_new_r2;
    reg [27:0] B_new_r2;

    reg [27:0] R_new_r3;
    reg [27:0] G_new_r3;
    reg [27:0] B_new_r3;

    reg [27:0] R_new_r4;
    reg [27:0] G_new_r4;
    reg [27:0] B_new_r4;


    wire   [7:0] rgb888_r_d1[0:3];
    wire   [7:0] rgb888_g_d1[0:3];
    wire   [7:0] rgb888_b_d1[0:3];

    assign  rgb888_r_d1[0] = data_d1[16+:8];
    assign  rgb888_g_d1[0] = data_d1[8+:8];
    assign  rgb888_b_d1[0] = data_d1[0+:8];

    assign  rgb888_r_d1[1] = data_d1[40+:8];
    assign  rgb888_g_d1[1] = data_d1[32+:8];
    assign  rgb888_b_d1[1] = data_d1[24+:8];

    assign  rgb888_r_d1[2] = data_d1[64+:8];
    assign  rgb888_g_d1[2] = data_d1[56+:8];
    assign  rgb888_b_d1[2] = data_d1[48+:8];

    assign  rgb888_r_d1[3] = data_d1[88+:8];
    assign  rgb888_g_d1[3] = data_d1[80+:8];
    assign  rgb888_b_d1[3] = data_d1[72+:8];
// �����µ�RGBֵ��Ӧ������
always @(posedge I_clk or negedge I_rst_n)begin 
    if(!I_rst_n)begin
        R_new_r1 <= 0;
        G_new_r1 <= 0;
        B_new_r1 <= 0;

        R_new_r2 <= 0;
        G_new_r2 <= 0;
        B_new_r2 <= 0;

        R_new_r3 <= 0;
        G_new_r3 <= 0;
        B_new_r3 <= 0;

        R_new_r4 <= 0;
        G_new_r4 <= 0;
        B_new_r4 <= 0;
    end
    else if(valid_d1) begin
        R_new_r1 <= in_r_r1 * rgb888_r_d1[0];
        G_new_r1 <=           rgb888_g_d1[0];
        B_new_r1 <= in_b_r1 * rgb888_b_d1[0];

        R_new_r2 <= in_r_r1 * rgb888_r_d1[1];
        G_new_r2 <=           rgb888_g_d1[1];
        B_new_r2 <= in_b_r1 * rgb888_b_d1[1];

        R_new_r3 <= in_r_r1 * rgb888_r_d1[2];
        G_new_r3 <=           rgb888_g_d1[2];
        B_new_r3 <= in_b_r1 * rgb888_b_d1[2];

        R_new_r4 <= in_r_r1 * rgb888_r_d1[3];
        G_new_r4 <=           rgb888_g_d1[3];
        B_new_r4 <= in_b_r1 * rgb888_b_d1[3];
    end
end

/*****************************************************************
                            ??????????                                      
*****************************************************************/

    wire [7:0] R_new_x1;
    wire [7:0] G_new_x1;
    wire [7:0] B_new_x1;

    wire [7:0] R_new_x2;
    wire [7:0] G_new_x2;
    wire [7:0] B_new_x2;

    wire [7:0] R_new_x3;
    wire [7:0] G_new_x3;
    wire [7:0] B_new_x3;

    wire [7:0] R_new_x4;
    wire [7:0] G_new_x4;
    wire [7:0] B_new_x4;

    assign R_new_x1 = (R_new_r1[27:24])?255:R_new_r1[23:16];
    assign G_new_x1 =  G_new_r1;
    assign B_new_x1 = (B_new_r1[27:24])?255:B_new_r1[23:16];

    assign R_new_x2 = (R_new_r2[27:24])?255:R_new_r2[23:16];
    assign G_new_x2 =  G_new_r2;
    assign B_new_x2 = (B_new_r2[27:24])?255:B_new_r2[23:16];

    assign R_new_x3 = (R_new_r3[27:24])?255:R_new_r3[23:16];
    assign G_new_x3 =  G_new_r3;
    assign B_new_x3 = (B_new_r3[27:24])?255:B_new_r3[23:16];

    assign R_new_x4 = (R_new_r4[27:24])?255:R_new_r4[23:16];
    assign G_new_x4 =  G_new_r4;
    assign B_new_x4 = (B_new_r4[27:24])?255:B_new_r4[23:16];
/*****************************************************************
                           ??????                                       
*****************************************************************/

    reg valid_d2,I_tuser_r2;
    always @(posedge I_clk or negedge I_rst_n) begin
        if(!I_rst_n)begin
            valid_d2 <= 0;
            I_tuser_r2 <= 0;
        end
        else begin
            valid_d2 <= valid_d1;
            I_tuser_r2 <= I_tuser_r1;
        end
    end


    assign  O_tlast  = (valid_d1 == 0) && (valid_d2 == 1);   
    assign  O_tuser  = I_tuser_r2 ;   
    assign  O_tvalid = valid_d2;

    assign  O_tdata = O_tvalid?{R_new_x4,G_new_x4,B_new_x4,
                       R_new_x3,G_new_x3,B_new_x3,
                       R_new_x2,G_new_x2,B_new_x2,
                       R_new_x1,G_new_x1,B_new_x1}:0;
    // assign O_t_data = {R_new[7-:5],G_new[7-:6],B_new[7-:5]};
    assign  I_tready = O_tready;
 
endmodule



